
	/* verilator lint_off COMBDLY */
	module rom_array_layer_2 #(
	parameter WIDTH=16,
	parameter KERNEL=1,
	parameter ADDR=8,
	parameter NUM=512)
	(
		input [ADDR-1:0] address ,
		output [WIDTH-1:0] rom_out [0:NUM-1]
	);	
	

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_1 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_2 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_3 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_4 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_5 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_6 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_7 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_8 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_9 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_10 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_11 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_12 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_13 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_14 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_15 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_16 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_17 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_18 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_19 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_20 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_21 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_22 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_23 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_24 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_25 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_26 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_27 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_28 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_29 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_30 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_31 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_32 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_33 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_34 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_35 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_36 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_37 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_38 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_39 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_40 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_41 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_42 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_43 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_44 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_45 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_46 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_47 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_48 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_49 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_50 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_51 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_52 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_53 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_54 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_55 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_56 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_57 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_58 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_59 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_60 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_61 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_62 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_63 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_64 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_65 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_66 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_67 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_68 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_69 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_70 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_71 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_72 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_73 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_74 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_75 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_76 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_77 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_78 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_79 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_80 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_81 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_82 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_83 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_84 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_85 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_86 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_87 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_88 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_89 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_90 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_91 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_92 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_93 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_94 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_95 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_96 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_97 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_98 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_99 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_100 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_101 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_102 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_103 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_104 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_105 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_106 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_107 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_108 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_109 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_110 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_111 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_112 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_113 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_114 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_115 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_116 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_117 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_118 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_119 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_120 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_121 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_122 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_123 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_124 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_125 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_126 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_127 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_128 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_129 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_130 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_131 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_132 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_133 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_134 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_135 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_136 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_137 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_138 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_139 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_140 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_141 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_142 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_143 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_144 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_145 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_146 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_147 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_148 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_149 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_150 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_151 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_152 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_153 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_154 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_155 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_156 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_157 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_158 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_159 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_160 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_161 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_162 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_163 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_164 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_165 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_166 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_167 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_168 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_169 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_170 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_171 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_172 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_173 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_174 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_175 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_176 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_177 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_178 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_179 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_180 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_181 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_182 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_183 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_184 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_185 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_186 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_187 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_188 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_189 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_190 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_191 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_192 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_193 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_194 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_195 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_196 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_197 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_198 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_199 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_200 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_201 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_202 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_203 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_204 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_205 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_206 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_207 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_208 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_209 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_210 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_211 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_212 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_213 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_214 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_215 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_216 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_217 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_218 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_219 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_220 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_221 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_222 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_223 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_224 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_225 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_226 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_227 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_228 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_229 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_230 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_231 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_232 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_233 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_234 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_235 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_236 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_237 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_238 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_239 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_240 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_241 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_242 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_243 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_244 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_245 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_246 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_247 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_248 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_249 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_250 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_251 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_252 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_253 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_254 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_255 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_256 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_257 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_258 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_259 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_260 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_261 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_262 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_263 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_264 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_265 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_266 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_267 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_268 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_269 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_270 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_271 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_272 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_273 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_274 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_275 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_276 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_277 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_278 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_279 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_280 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_281 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_282 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_283 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_284 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_285 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_286 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_287 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_288 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_289 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_290 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_291 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_292 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_293 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_294 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_295 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_296 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_297 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_298 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_299 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_300 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_301 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_302 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_303 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_304 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_305 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_306 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_307 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_308 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_309 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_310 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_311 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_312 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_313 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_314 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_315 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_316 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_317 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_318 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_319 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_320 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_321 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_322 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_323 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_324 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_325 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_326 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_327 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_328 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_329 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_330 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_331 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_332 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_333 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_334 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_335 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_336 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_337 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_338 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_339 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_340 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_341 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_342 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_343 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_344 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_345 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_346 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_347 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_348 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_349 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_350 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_351 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_352 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_353 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_354 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_355 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_356 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_357 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_358 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_359 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_360 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_361 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_362 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_363 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_364 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_365 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_366 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_367 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_368 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_369 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_370 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_371 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_372 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_373 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_374 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_375 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_376 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_377 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_378 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_379 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_380 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_381 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_382 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_383 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_384 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_385 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_386 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_387 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_388 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_389 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_390 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_391 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_392 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_393 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_394 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_395 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_396 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_397 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_398 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_399 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_400 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_401 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_402 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_403 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_404 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_405 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_406 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_407 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_408 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_409 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_410 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_411 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_412 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_413 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_414 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_415 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_416 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_417 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_418 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_419 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_420 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_421 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_422 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_423 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_424 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_425 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_426 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_427 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_428 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_429 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_430 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_431 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_432 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_433 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_434 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_435 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_436 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_437 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_438 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_439 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_440 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_441 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_442 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_443 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_444 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_445 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_446 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_447 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_448 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_449 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_450 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_451 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_452 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_453 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_454 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_455 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_456 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_457 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_458 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_459 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_460 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_461 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_462 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_463 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_464 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_465 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_466 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_467 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_468 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_469 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_470 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_471 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_472 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_473 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_474 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_475 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_476 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_477 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_478 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_479 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_480 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_481 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_482 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_483 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_484 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_485 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_486 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_487 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_488 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_489 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_490 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_491 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_492 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_493 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_494 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_495 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_496 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_497 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_498 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_499 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_500 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_501 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_502 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_503 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_504 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_505 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_506 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_507 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_508 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_509 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_510 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_511 [0:2**ADDR-1] ;

  	(* rom_style="{distributed}" *)
	reg [WIDTH-1:0] rom_512 [0:2**ADDR-1] ;
initial begin
$readmemb("extend_file_1.mem",rom_1,0,2**ADDR-1);
$readmemb("extend_file_2.mem",rom_2,0,2**ADDR-1);
$readmemb("extend_file_3.mem",rom_3,0,2**ADDR-1);
$readmemb("extend_file_4.mem",rom_4,0,2**ADDR-1);
$readmemb("extend_file_5.mem",rom_5,0,2**ADDR-1);
$readmemb("extend_file_6.mem",rom_6,0,2**ADDR-1);
$readmemb("extend_file_7.mem",rom_7,0,2**ADDR-1);
$readmemb("extend_file_8.mem",rom_8,0,2**ADDR-1);
$readmemb("extend_file_9.mem",rom_9,0,2**ADDR-1);
$readmemb("extend_file_10.mem",rom_10,0,2**ADDR-1);
$readmemb("extend_file_11.mem",rom_11,0,2**ADDR-1);
$readmemb("extend_file_12.mem",rom_12,0,2**ADDR-1);
$readmemb("extend_file_13.mem",rom_13,0,2**ADDR-1);
$readmemb("extend_file_14.mem",rom_14,0,2**ADDR-1);
$readmemb("extend_file_15.mem",rom_15,0,2**ADDR-1);
$readmemb("extend_file_16.mem",rom_16,0,2**ADDR-1);
$readmemb("extend_file_17.mem",rom_17,0,2**ADDR-1);
$readmemb("extend_file_18.mem",rom_18,0,2**ADDR-1);
$readmemb("extend_file_19.mem",rom_19,0,2**ADDR-1);
$readmemb("extend_file_20.mem",rom_20,0,2**ADDR-1);
$readmemb("extend_file_21.mem",rom_21,0,2**ADDR-1);
$readmemb("extend_file_22.mem",rom_22,0,2**ADDR-1);
$readmemb("extend_file_23.mem",rom_23,0,2**ADDR-1);
$readmemb("extend_file_24.mem",rom_24,0,2**ADDR-1);
$readmemb("extend_file_25.mem",rom_25,0,2**ADDR-1);
$readmemb("extend_file_26.mem",rom_26,0,2**ADDR-1);
$readmemb("extend_file_27.mem",rom_27,0,2**ADDR-1);
$readmemb("extend_file_28.mem",rom_28,0,2**ADDR-1);
$readmemb("extend_file_29.mem",rom_29,0,2**ADDR-1);
$readmemb("extend_file_30.mem",rom_30,0,2**ADDR-1);
$readmemb("extend_file_31.mem",rom_31,0,2**ADDR-1);
$readmemb("extend_file_32.mem",rom_32,0,2**ADDR-1);
$readmemb("extend_file_33.mem",rom_33,0,2**ADDR-1);
$readmemb("extend_file_34.mem",rom_34,0,2**ADDR-1);
$readmemb("extend_file_35.mem",rom_35,0,2**ADDR-1);
$readmemb("extend_file_36.mem",rom_36,0,2**ADDR-1);
$readmemb("extend_file_37.mem",rom_37,0,2**ADDR-1);
$readmemb("extend_file_38.mem",rom_38,0,2**ADDR-1);
$readmemb("extend_file_39.mem",rom_39,0,2**ADDR-1);
$readmemb("extend_file_40.mem",rom_40,0,2**ADDR-1);
$readmemb("extend_file_41.mem",rom_41,0,2**ADDR-1);
$readmemb("extend_file_42.mem",rom_42,0,2**ADDR-1);
$readmemb("extend_file_43.mem",rom_43,0,2**ADDR-1);
$readmemb("extend_file_44.mem",rom_44,0,2**ADDR-1);
$readmemb("extend_file_45.mem",rom_45,0,2**ADDR-1);
$readmemb("extend_file_46.mem",rom_46,0,2**ADDR-1);
$readmemb("extend_file_47.mem",rom_47,0,2**ADDR-1);
$readmemb("extend_file_48.mem",rom_48,0,2**ADDR-1);
$readmemb("extend_file_49.mem",rom_49,0,2**ADDR-1);
$readmemb("extend_file_50.mem",rom_50,0,2**ADDR-1);
$readmemb("extend_file_51.mem",rom_51,0,2**ADDR-1);
$readmemb("extend_file_52.mem",rom_52,0,2**ADDR-1);
$readmemb("extend_file_53.mem",rom_53,0,2**ADDR-1);
$readmemb("extend_file_54.mem",rom_54,0,2**ADDR-1);
$readmemb("extend_file_55.mem",rom_55,0,2**ADDR-1);
$readmemb("extend_file_56.mem",rom_56,0,2**ADDR-1);
$readmemb("extend_file_57.mem",rom_57,0,2**ADDR-1);
$readmemb("extend_file_58.mem",rom_58,0,2**ADDR-1);
$readmemb("extend_file_59.mem",rom_59,0,2**ADDR-1);
$readmemb("extend_file_60.mem",rom_60,0,2**ADDR-1);
$readmemb("extend_file_61.mem",rom_61,0,2**ADDR-1);
$readmemb("extend_file_62.mem",rom_62,0,2**ADDR-1);
$readmemb("extend_file_63.mem",rom_63,0,2**ADDR-1);
$readmemb("extend_file_64.mem",rom_64,0,2**ADDR-1);
$readmemb("extend_file_65.mem",rom_65,0,2**ADDR-1);
$readmemb("extend_file_66.mem",rom_66,0,2**ADDR-1);
$readmemb("extend_file_67.mem",rom_67,0,2**ADDR-1);
$readmemb("extend_file_68.mem",rom_68,0,2**ADDR-1);
$readmemb("extend_file_69.mem",rom_69,0,2**ADDR-1);
$readmemb("extend_file_70.mem",rom_70,0,2**ADDR-1);
$readmemb("extend_file_71.mem",rom_71,0,2**ADDR-1);
$readmemb("extend_file_72.mem",rom_72,0,2**ADDR-1);
$readmemb("extend_file_73.mem",rom_73,0,2**ADDR-1);
$readmemb("extend_file_74.mem",rom_74,0,2**ADDR-1);
$readmemb("extend_file_75.mem",rom_75,0,2**ADDR-1);
$readmemb("extend_file_76.mem",rom_76,0,2**ADDR-1);
$readmemb("extend_file_77.mem",rom_77,0,2**ADDR-1);
$readmemb("extend_file_78.mem",rom_78,0,2**ADDR-1);
$readmemb("extend_file_79.mem",rom_79,0,2**ADDR-1);
$readmemb("extend_file_80.mem",rom_80,0,2**ADDR-1);
$readmemb("extend_file_81.mem",rom_81,0,2**ADDR-1);
$readmemb("extend_file_82.mem",rom_82,0,2**ADDR-1);
$readmemb("extend_file_83.mem",rom_83,0,2**ADDR-1);
$readmemb("extend_file_84.mem",rom_84,0,2**ADDR-1);
$readmemb("extend_file_85.mem",rom_85,0,2**ADDR-1);
$readmemb("extend_file_86.mem",rom_86,0,2**ADDR-1);
$readmemb("extend_file_87.mem",rom_87,0,2**ADDR-1);
$readmemb("extend_file_88.mem",rom_88,0,2**ADDR-1);
$readmemb("extend_file_89.mem",rom_89,0,2**ADDR-1);
$readmemb("extend_file_90.mem",rom_90,0,2**ADDR-1);
$readmemb("extend_file_91.mem",rom_91,0,2**ADDR-1);
$readmemb("extend_file_92.mem",rom_92,0,2**ADDR-1);
$readmemb("extend_file_93.mem",rom_93,0,2**ADDR-1);
$readmemb("extend_file_94.mem",rom_94,0,2**ADDR-1);
$readmemb("extend_file_95.mem",rom_95,0,2**ADDR-1);
$readmemb("extend_file_96.mem",rom_96,0,2**ADDR-1);
$readmemb("extend_file_97.mem",rom_97,0,2**ADDR-1);
$readmemb("extend_file_98.mem",rom_98,0,2**ADDR-1);
$readmemb("extend_file_99.mem",rom_99,0,2**ADDR-1);
$readmemb("extend_file_100.mem",rom_100,0,2**ADDR-1);
$readmemb("extend_file_101.mem",rom_101,0,2**ADDR-1);
$readmemb("extend_file_102.mem",rom_102,0,2**ADDR-1);
$readmemb("extend_file_103.mem",rom_103,0,2**ADDR-1);
$readmemb("extend_file_104.mem",rom_104,0,2**ADDR-1);
$readmemb("extend_file_105.mem",rom_105,0,2**ADDR-1);
$readmemb("extend_file_106.mem",rom_106,0,2**ADDR-1);
$readmemb("extend_file_107.mem",rom_107,0,2**ADDR-1);
$readmemb("extend_file_108.mem",rom_108,0,2**ADDR-1);
$readmemb("extend_file_109.mem",rom_109,0,2**ADDR-1);
$readmemb("extend_file_110.mem",rom_110,0,2**ADDR-1);
$readmemb("extend_file_111.mem",rom_111,0,2**ADDR-1);
$readmemb("extend_file_112.mem",rom_112,0,2**ADDR-1);
$readmemb("extend_file_113.mem",rom_113,0,2**ADDR-1);
$readmemb("extend_file_114.mem",rom_114,0,2**ADDR-1);
$readmemb("extend_file_115.mem",rom_115,0,2**ADDR-1);
$readmemb("extend_file_116.mem",rom_116,0,2**ADDR-1);
$readmemb("extend_file_117.mem",rom_117,0,2**ADDR-1);
$readmemb("extend_file_118.mem",rom_118,0,2**ADDR-1);
$readmemb("extend_file_119.mem",rom_119,0,2**ADDR-1);
$readmemb("extend_file_120.mem",rom_120,0,2**ADDR-1);
$readmemb("extend_file_121.mem",rom_121,0,2**ADDR-1);
$readmemb("extend_file_122.mem",rom_122,0,2**ADDR-1);
$readmemb("extend_file_123.mem",rom_123,0,2**ADDR-1);
$readmemb("extend_file_124.mem",rom_124,0,2**ADDR-1);
$readmemb("extend_file_125.mem",rom_125,0,2**ADDR-1);
$readmemb("extend_file_126.mem",rom_126,0,2**ADDR-1);
$readmemb("extend_file_127.mem",rom_127,0,2**ADDR-1);
$readmemb("extend_file_128.mem",rom_128,0,2**ADDR-1);
$readmemb("extend_file_129.mem",rom_129,0,2**ADDR-1);
$readmemb("extend_file_130.mem",rom_130,0,2**ADDR-1);
$readmemb("extend_file_131.mem",rom_131,0,2**ADDR-1);
$readmemb("extend_file_132.mem",rom_132,0,2**ADDR-1);
$readmemb("extend_file_133.mem",rom_133,0,2**ADDR-1);
$readmemb("extend_file_134.mem",rom_134,0,2**ADDR-1);
$readmemb("extend_file_135.mem",rom_135,0,2**ADDR-1);
$readmemb("extend_file_136.mem",rom_136,0,2**ADDR-1);
$readmemb("extend_file_137.mem",rom_137,0,2**ADDR-1);
$readmemb("extend_file_138.mem",rom_138,0,2**ADDR-1);
$readmemb("extend_file_139.mem",rom_139,0,2**ADDR-1);
$readmemb("extend_file_140.mem",rom_140,0,2**ADDR-1);
$readmemb("extend_file_141.mem",rom_141,0,2**ADDR-1);
$readmemb("extend_file_142.mem",rom_142,0,2**ADDR-1);
$readmemb("extend_file_143.mem",rom_143,0,2**ADDR-1);
$readmemb("extend_file_144.mem",rom_144,0,2**ADDR-1);
$readmemb("extend_file_145.mem",rom_145,0,2**ADDR-1);
$readmemb("extend_file_146.mem",rom_146,0,2**ADDR-1);
$readmemb("extend_file_147.mem",rom_147,0,2**ADDR-1);
$readmemb("extend_file_148.mem",rom_148,0,2**ADDR-1);
$readmemb("extend_file_149.mem",rom_149,0,2**ADDR-1);
$readmemb("extend_file_150.mem",rom_150,0,2**ADDR-1);
$readmemb("extend_file_151.mem",rom_151,0,2**ADDR-1);
$readmemb("extend_file_152.mem",rom_152,0,2**ADDR-1);
$readmemb("extend_file_153.mem",rom_153,0,2**ADDR-1);
$readmemb("extend_file_154.mem",rom_154,0,2**ADDR-1);
$readmemb("extend_file_155.mem",rom_155,0,2**ADDR-1);
$readmemb("extend_file_156.mem",rom_156,0,2**ADDR-1);
$readmemb("extend_file_157.mem",rom_157,0,2**ADDR-1);
$readmemb("extend_file_158.mem",rom_158,0,2**ADDR-1);
$readmemb("extend_file_159.mem",rom_159,0,2**ADDR-1);
$readmemb("extend_file_160.mem",rom_160,0,2**ADDR-1);
$readmemb("extend_file_161.mem",rom_161,0,2**ADDR-1);
$readmemb("extend_file_162.mem",rom_162,0,2**ADDR-1);
$readmemb("extend_file_163.mem",rom_163,0,2**ADDR-1);
$readmemb("extend_file_164.mem",rom_164,0,2**ADDR-1);
$readmemb("extend_file_165.mem",rom_165,0,2**ADDR-1);
$readmemb("extend_file_166.mem",rom_166,0,2**ADDR-1);
$readmemb("extend_file_167.mem",rom_167,0,2**ADDR-1);
$readmemb("extend_file_168.mem",rom_168,0,2**ADDR-1);
$readmemb("extend_file_169.mem",rom_169,0,2**ADDR-1);
$readmemb("extend_file_170.mem",rom_170,0,2**ADDR-1);
$readmemb("extend_file_171.mem",rom_171,0,2**ADDR-1);
$readmemb("extend_file_172.mem",rom_172,0,2**ADDR-1);
$readmemb("extend_file_173.mem",rom_173,0,2**ADDR-1);
$readmemb("extend_file_174.mem",rom_174,0,2**ADDR-1);
$readmemb("extend_file_175.mem",rom_175,0,2**ADDR-1);
$readmemb("extend_file_176.mem",rom_176,0,2**ADDR-1);
$readmemb("extend_file_177.mem",rom_177,0,2**ADDR-1);
$readmemb("extend_file_178.mem",rom_178,0,2**ADDR-1);
$readmemb("extend_file_179.mem",rom_179,0,2**ADDR-1);
$readmemb("extend_file_180.mem",rom_180,0,2**ADDR-1);
$readmemb("extend_file_181.mem",rom_181,0,2**ADDR-1);
$readmemb("extend_file_182.mem",rom_182,0,2**ADDR-1);
$readmemb("extend_file_183.mem",rom_183,0,2**ADDR-1);
$readmemb("extend_file_184.mem",rom_184,0,2**ADDR-1);
$readmemb("extend_file_185.mem",rom_185,0,2**ADDR-1);
$readmemb("extend_file_186.mem",rom_186,0,2**ADDR-1);
$readmemb("extend_file_187.mem",rom_187,0,2**ADDR-1);
$readmemb("extend_file_188.mem",rom_188,0,2**ADDR-1);
$readmemb("extend_file_189.mem",rom_189,0,2**ADDR-1);
$readmemb("extend_file_190.mem",rom_190,0,2**ADDR-1);
$readmemb("extend_file_191.mem",rom_191,0,2**ADDR-1);
$readmemb("extend_file_192.mem",rom_192,0,2**ADDR-1);
$readmemb("extend_file_193.mem",rom_193,0,2**ADDR-1);
$readmemb("extend_file_194.mem",rom_194,0,2**ADDR-1);
$readmemb("extend_file_195.mem",rom_195,0,2**ADDR-1);
$readmemb("extend_file_196.mem",rom_196,0,2**ADDR-1);
$readmemb("extend_file_197.mem",rom_197,0,2**ADDR-1);
$readmemb("extend_file_198.mem",rom_198,0,2**ADDR-1);
$readmemb("extend_file_199.mem",rom_199,0,2**ADDR-1);
$readmemb("extend_file_200.mem",rom_200,0,2**ADDR-1);
$readmemb("extend_file_201.mem",rom_201,0,2**ADDR-1);
$readmemb("extend_file_202.mem",rom_202,0,2**ADDR-1);
$readmemb("extend_file_203.mem",rom_203,0,2**ADDR-1);
$readmemb("extend_file_204.mem",rom_204,0,2**ADDR-1);
$readmemb("extend_file_205.mem",rom_205,0,2**ADDR-1);
$readmemb("extend_file_206.mem",rom_206,0,2**ADDR-1);
$readmemb("extend_file_207.mem",rom_207,0,2**ADDR-1);
$readmemb("extend_file_208.mem",rom_208,0,2**ADDR-1);
$readmemb("extend_file_209.mem",rom_209,0,2**ADDR-1);
$readmemb("extend_file_210.mem",rom_210,0,2**ADDR-1);
$readmemb("extend_file_211.mem",rom_211,0,2**ADDR-1);
$readmemb("extend_file_212.mem",rom_212,0,2**ADDR-1);
$readmemb("extend_file_213.mem",rom_213,0,2**ADDR-1);
$readmemb("extend_file_214.mem",rom_214,0,2**ADDR-1);
$readmemb("extend_file_215.mem",rom_215,0,2**ADDR-1);
$readmemb("extend_file_216.mem",rom_216,0,2**ADDR-1);
$readmemb("extend_file_217.mem",rom_217,0,2**ADDR-1);
$readmemb("extend_file_218.mem",rom_218,0,2**ADDR-1);
$readmemb("extend_file_219.mem",rom_219,0,2**ADDR-1);
$readmemb("extend_file_220.mem",rom_220,0,2**ADDR-1);
$readmemb("extend_file_221.mem",rom_221,0,2**ADDR-1);
$readmemb("extend_file_222.mem",rom_222,0,2**ADDR-1);
$readmemb("extend_file_223.mem",rom_223,0,2**ADDR-1);
$readmemb("extend_file_224.mem",rom_224,0,2**ADDR-1);
$readmemb("extend_file_225.mem",rom_225,0,2**ADDR-1);
$readmemb("extend_file_226.mem",rom_226,0,2**ADDR-1);
$readmemb("extend_file_227.mem",rom_227,0,2**ADDR-1);
$readmemb("extend_file_228.mem",rom_228,0,2**ADDR-1);
$readmemb("extend_file_229.mem",rom_229,0,2**ADDR-1);
$readmemb("extend_file_230.mem",rom_230,0,2**ADDR-1);
$readmemb("extend_file_231.mem",rom_231,0,2**ADDR-1);
$readmemb("extend_file_232.mem",rom_232,0,2**ADDR-1);
$readmemb("extend_file_233.mem",rom_233,0,2**ADDR-1);
$readmemb("extend_file_234.mem",rom_234,0,2**ADDR-1);
$readmemb("extend_file_235.mem",rom_235,0,2**ADDR-1);
$readmemb("extend_file_236.mem",rom_236,0,2**ADDR-1);
$readmemb("extend_file_237.mem",rom_237,0,2**ADDR-1);
$readmemb("extend_file_238.mem",rom_238,0,2**ADDR-1);
$readmemb("extend_file_239.mem",rom_239,0,2**ADDR-1);
$readmemb("extend_file_240.mem",rom_240,0,2**ADDR-1);
$readmemb("extend_file_241.mem",rom_241,0,2**ADDR-1);
$readmemb("extend_file_242.mem",rom_242,0,2**ADDR-1);
$readmemb("extend_file_243.mem",rom_243,0,2**ADDR-1);
$readmemb("extend_file_244.mem",rom_244,0,2**ADDR-1);
$readmemb("extend_file_245.mem",rom_245,0,2**ADDR-1);
$readmemb("extend_file_246.mem",rom_246,0,2**ADDR-1);
$readmemb("extend_file_247.mem",rom_247,0,2**ADDR-1);
$readmemb("extend_file_248.mem",rom_248,0,2**ADDR-1);
$readmemb("extend_file_249.mem",rom_249,0,2**ADDR-1);
$readmemb("extend_file_250.mem",rom_250,0,2**ADDR-1);
$readmemb("extend_file_251.mem",rom_251,0,2**ADDR-1);
$readmemb("extend_file_252.mem",rom_252,0,2**ADDR-1);
$readmemb("extend_file_253.mem",rom_253,0,2**ADDR-1);
$readmemb("extend_file_254.mem",rom_254,0,2**ADDR-1);
$readmemb("extend_file_255.mem",rom_255,0,2**ADDR-1);
$readmemb("extend_file_256.mem",rom_256,0,2**ADDR-1);
$readmemb("extend_file_257.mem",rom_257,0,2**ADDR-1);
$readmemb("extend_file_258.mem",rom_258,0,2**ADDR-1);
$readmemb("extend_file_259.mem",rom_259,0,2**ADDR-1);
$readmemb("extend_file_260.mem",rom_260,0,2**ADDR-1);
$readmemb("extend_file_261.mem",rom_261,0,2**ADDR-1);
$readmemb("extend_file_262.mem",rom_262,0,2**ADDR-1);
$readmemb("extend_file_263.mem",rom_263,0,2**ADDR-1);
$readmemb("extend_file_264.mem",rom_264,0,2**ADDR-1);
$readmemb("extend_file_265.mem",rom_265,0,2**ADDR-1);
$readmemb("extend_file_266.mem",rom_266,0,2**ADDR-1);
$readmemb("extend_file_267.mem",rom_267,0,2**ADDR-1);
$readmemb("extend_file_268.mem",rom_268,0,2**ADDR-1);
$readmemb("extend_file_269.mem",rom_269,0,2**ADDR-1);
$readmemb("extend_file_270.mem",rom_270,0,2**ADDR-1);
$readmemb("extend_file_271.mem",rom_271,0,2**ADDR-1);
$readmemb("extend_file_272.mem",rom_272,0,2**ADDR-1);
$readmemb("extend_file_273.mem",rom_273,0,2**ADDR-1);
$readmemb("extend_file_274.mem",rom_274,0,2**ADDR-1);
$readmemb("extend_file_275.mem",rom_275,0,2**ADDR-1);
$readmemb("extend_file_276.mem",rom_276,0,2**ADDR-1);
$readmemb("extend_file_277.mem",rom_277,0,2**ADDR-1);
$readmemb("extend_file_278.mem",rom_278,0,2**ADDR-1);
$readmemb("extend_file_279.mem",rom_279,0,2**ADDR-1);
$readmemb("extend_file_280.mem",rom_280,0,2**ADDR-1);
$readmemb("extend_file_281.mem",rom_281,0,2**ADDR-1);
$readmemb("extend_file_282.mem",rom_282,0,2**ADDR-1);
$readmemb("extend_file_283.mem",rom_283,0,2**ADDR-1);
$readmemb("extend_file_284.mem",rom_284,0,2**ADDR-1);
$readmemb("extend_file_285.mem",rom_285,0,2**ADDR-1);
$readmemb("extend_file_286.mem",rom_286,0,2**ADDR-1);
$readmemb("extend_file_287.mem",rom_287,0,2**ADDR-1);
$readmemb("extend_file_288.mem",rom_288,0,2**ADDR-1);
$readmemb("extend_file_289.mem",rom_289,0,2**ADDR-1);
$readmemb("extend_file_290.mem",rom_290,0,2**ADDR-1);
$readmemb("extend_file_291.mem",rom_291,0,2**ADDR-1);
$readmemb("extend_file_292.mem",rom_292,0,2**ADDR-1);
$readmemb("extend_file_293.mem",rom_293,0,2**ADDR-1);
$readmemb("extend_file_294.mem",rom_294,0,2**ADDR-1);
$readmemb("extend_file_295.mem",rom_295,0,2**ADDR-1);
$readmemb("extend_file_296.mem",rom_296,0,2**ADDR-1);
$readmemb("extend_file_297.mem",rom_297,0,2**ADDR-1);
$readmemb("extend_file_298.mem",rom_298,0,2**ADDR-1);
$readmemb("extend_file_299.mem",rom_299,0,2**ADDR-1);
$readmemb("extend_file_300.mem",rom_300,0,2**ADDR-1);
$readmemb("extend_file_301.mem",rom_301,0,2**ADDR-1);
$readmemb("extend_file_302.mem",rom_302,0,2**ADDR-1);
$readmemb("extend_file_303.mem",rom_303,0,2**ADDR-1);
$readmemb("extend_file_304.mem",rom_304,0,2**ADDR-1);
$readmemb("extend_file_305.mem",rom_305,0,2**ADDR-1);
$readmemb("extend_file_306.mem",rom_306,0,2**ADDR-1);
$readmemb("extend_file_307.mem",rom_307,0,2**ADDR-1);
$readmemb("extend_file_308.mem",rom_308,0,2**ADDR-1);
$readmemb("extend_file_309.mem",rom_309,0,2**ADDR-1);
$readmemb("extend_file_310.mem",rom_310,0,2**ADDR-1);
$readmemb("extend_file_311.mem",rom_311,0,2**ADDR-1);
$readmemb("extend_file_312.mem",rom_312,0,2**ADDR-1);
$readmemb("extend_file_313.mem",rom_313,0,2**ADDR-1);
$readmemb("extend_file_314.mem",rom_314,0,2**ADDR-1);
$readmemb("extend_file_315.mem",rom_315,0,2**ADDR-1);
$readmemb("extend_file_316.mem",rom_316,0,2**ADDR-1);
$readmemb("extend_file_317.mem",rom_317,0,2**ADDR-1);
$readmemb("extend_file_318.mem",rom_318,0,2**ADDR-1);
$readmemb("extend_file_319.mem",rom_319,0,2**ADDR-1);
$readmemb("extend_file_320.mem",rom_320,0,2**ADDR-1);
$readmemb("extend_file_321.mem",rom_321,0,2**ADDR-1);
$readmemb("extend_file_322.mem",rom_322,0,2**ADDR-1);
$readmemb("extend_file_323.mem",rom_323,0,2**ADDR-1);
$readmemb("extend_file_324.mem",rom_324,0,2**ADDR-1);
$readmemb("extend_file_325.mem",rom_325,0,2**ADDR-1);
$readmemb("extend_file_326.mem",rom_326,0,2**ADDR-1);
$readmemb("extend_file_327.mem",rom_327,0,2**ADDR-1);
$readmemb("extend_file_328.mem",rom_328,0,2**ADDR-1);
$readmemb("extend_file_329.mem",rom_329,0,2**ADDR-1);
$readmemb("extend_file_330.mem",rom_330,0,2**ADDR-1);
$readmemb("extend_file_331.mem",rom_331,0,2**ADDR-1);
$readmemb("extend_file_332.mem",rom_332,0,2**ADDR-1);
$readmemb("extend_file_333.mem",rom_333,0,2**ADDR-1);
$readmemb("extend_file_334.mem",rom_334,0,2**ADDR-1);
$readmemb("extend_file_335.mem",rom_335,0,2**ADDR-1);
$readmemb("extend_file_336.mem",rom_336,0,2**ADDR-1);
$readmemb("extend_file_337.mem",rom_337,0,2**ADDR-1);
$readmemb("extend_file_338.mem",rom_338,0,2**ADDR-1);
$readmemb("extend_file_339.mem",rom_339,0,2**ADDR-1);
$readmemb("extend_file_340.mem",rom_340,0,2**ADDR-1);
$readmemb("extend_file_341.mem",rom_341,0,2**ADDR-1);
$readmemb("extend_file_342.mem",rom_342,0,2**ADDR-1);
$readmemb("extend_file_343.mem",rom_343,0,2**ADDR-1);
$readmemb("extend_file_344.mem",rom_344,0,2**ADDR-1);
$readmemb("extend_file_345.mem",rom_345,0,2**ADDR-1);
$readmemb("extend_file_346.mem",rom_346,0,2**ADDR-1);
$readmemb("extend_file_347.mem",rom_347,0,2**ADDR-1);
$readmemb("extend_file_348.mem",rom_348,0,2**ADDR-1);
$readmemb("extend_file_349.mem",rom_349,0,2**ADDR-1);
$readmemb("extend_file_350.mem",rom_350,0,2**ADDR-1);
$readmemb("extend_file_351.mem",rom_351,0,2**ADDR-1);
$readmemb("extend_file_352.mem",rom_352,0,2**ADDR-1);
$readmemb("extend_file_353.mem",rom_353,0,2**ADDR-1);
$readmemb("extend_file_354.mem",rom_354,0,2**ADDR-1);
$readmemb("extend_file_355.mem",rom_355,0,2**ADDR-1);
$readmemb("extend_file_356.mem",rom_356,0,2**ADDR-1);
$readmemb("extend_file_357.mem",rom_357,0,2**ADDR-1);
$readmemb("extend_file_358.mem",rom_358,0,2**ADDR-1);
$readmemb("extend_file_359.mem",rom_359,0,2**ADDR-1);
$readmemb("extend_file_360.mem",rom_360,0,2**ADDR-1);
$readmemb("extend_file_361.mem",rom_361,0,2**ADDR-1);
$readmemb("extend_file_362.mem",rom_362,0,2**ADDR-1);
$readmemb("extend_file_363.mem",rom_363,0,2**ADDR-1);
$readmemb("extend_file_364.mem",rom_364,0,2**ADDR-1);
$readmemb("extend_file_365.mem",rom_365,0,2**ADDR-1);
$readmemb("extend_file_366.mem",rom_366,0,2**ADDR-1);
$readmemb("extend_file_367.mem",rom_367,0,2**ADDR-1);
$readmemb("extend_file_368.mem",rom_368,0,2**ADDR-1);
$readmemb("extend_file_369.mem",rom_369,0,2**ADDR-1);
$readmemb("extend_file_370.mem",rom_370,0,2**ADDR-1);
$readmemb("extend_file_371.mem",rom_371,0,2**ADDR-1);
$readmemb("extend_file_372.mem",rom_372,0,2**ADDR-1);
$readmemb("extend_file_373.mem",rom_373,0,2**ADDR-1);
$readmemb("extend_file_374.mem",rom_374,0,2**ADDR-1);
$readmemb("extend_file_375.mem",rom_375,0,2**ADDR-1);
$readmemb("extend_file_376.mem",rom_376,0,2**ADDR-1);
$readmemb("extend_file_377.mem",rom_377,0,2**ADDR-1);
$readmemb("extend_file_378.mem",rom_378,0,2**ADDR-1);
$readmemb("extend_file_379.mem",rom_379,0,2**ADDR-1);
$readmemb("extend_file_380.mem",rom_380,0,2**ADDR-1);
$readmemb("extend_file_381.mem",rom_381,0,2**ADDR-1);
$readmemb("extend_file_382.mem",rom_382,0,2**ADDR-1);
$readmemb("extend_file_383.mem",rom_383,0,2**ADDR-1);
$readmemb("extend_file_384.mem",rom_384,0,2**ADDR-1);
$readmemb("extend_file_385.mem",rom_385,0,2**ADDR-1);
$readmemb("extend_file_386.mem",rom_386,0,2**ADDR-1);
$readmemb("extend_file_387.mem",rom_387,0,2**ADDR-1);
$readmemb("extend_file_388.mem",rom_388,0,2**ADDR-1);
$readmemb("extend_file_389.mem",rom_389,0,2**ADDR-1);
$readmemb("extend_file_390.mem",rom_390,0,2**ADDR-1);
$readmemb("extend_file_391.mem",rom_391,0,2**ADDR-1);
$readmemb("extend_file_392.mem",rom_392,0,2**ADDR-1);
$readmemb("extend_file_393.mem",rom_393,0,2**ADDR-1);
$readmemb("extend_file_394.mem",rom_394,0,2**ADDR-1);
$readmemb("extend_file_395.mem",rom_395,0,2**ADDR-1);
$readmemb("extend_file_396.mem",rom_396,0,2**ADDR-1);
$readmemb("extend_file_397.mem",rom_397,0,2**ADDR-1);
$readmemb("extend_file_398.mem",rom_398,0,2**ADDR-1);
$readmemb("extend_file_399.mem",rom_399,0,2**ADDR-1);
$readmemb("extend_file_400.mem",rom_400,0,2**ADDR-1);
$readmemb("extend_file_401.mem",rom_401,0,2**ADDR-1);
$readmemb("extend_file_402.mem",rom_402,0,2**ADDR-1);
$readmemb("extend_file_403.mem",rom_403,0,2**ADDR-1);
$readmemb("extend_file_404.mem",rom_404,0,2**ADDR-1);
$readmemb("extend_file_405.mem",rom_405,0,2**ADDR-1);
$readmemb("extend_file_406.mem",rom_406,0,2**ADDR-1);
$readmemb("extend_file_407.mem",rom_407,0,2**ADDR-1);
$readmemb("extend_file_408.mem",rom_408,0,2**ADDR-1);
$readmemb("extend_file_409.mem",rom_409,0,2**ADDR-1);
$readmemb("extend_file_410.mem",rom_410,0,2**ADDR-1);
$readmemb("extend_file_411.mem",rom_411,0,2**ADDR-1);
$readmemb("extend_file_412.mem",rom_412,0,2**ADDR-1);
$readmemb("extend_file_413.mem",rom_413,0,2**ADDR-1);
$readmemb("extend_file_414.mem",rom_414,0,2**ADDR-1);
$readmemb("extend_file_415.mem",rom_415,0,2**ADDR-1);
$readmemb("extend_file_416.mem",rom_416,0,2**ADDR-1);
$readmemb("extend_file_417.mem",rom_417,0,2**ADDR-1);
$readmemb("extend_file_418.mem",rom_418,0,2**ADDR-1);
$readmemb("extend_file_419.mem",rom_419,0,2**ADDR-1);
$readmemb("extend_file_420.mem",rom_420,0,2**ADDR-1);
$readmemb("extend_file_421.mem",rom_421,0,2**ADDR-1);
$readmemb("extend_file_422.mem",rom_422,0,2**ADDR-1);
$readmemb("extend_file_423.mem",rom_423,0,2**ADDR-1);
$readmemb("extend_file_424.mem",rom_424,0,2**ADDR-1);
$readmemb("extend_file_425.mem",rom_425,0,2**ADDR-1);
$readmemb("extend_file_426.mem",rom_426,0,2**ADDR-1);
$readmemb("extend_file_427.mem",rom_427,0,2**ADDR-1);
$readmemb("extend_file_428.mem",rom_428,0,2**ADDR-1);
$readmemb("extend_file_429.mem",rom_429,0,2**ADDR-1);
$readmemb("extend_file_430.mem",rom_430,0,2**ADDR-1);
$readmemb("extend_file_431.mem",rom_431,0,2**ADDR-1);
$readmemb("extend_file_432.mem",rom_432,0,2**ADDR-1);
$readmemb("extend_file_433.mem",rom_433,0,2**ADDR-1);
$readmemb("extend_file_434.mem",rom_434,0,2**ADDR-1);
$readmemb("extend_file_435.mem",rom_435,0,2**ADDR-1);
$readmemb("extend_file_436.mem",rom_436,0,2**ADDR-1);
$readmemb("extend_file_437.mem",rom_437,0,2**ADDR-1);
$readmemb("extend_file_438.mem",rom_438,0,2**ADDR-1);
$readmemb("extend_file_439.mem",rom_439,0,2**ADDR-1);
$readmemb("extend_file_440.mem",rom_440,0,2**ADDR-1);
$readmemb("extend_file_441.mem",rom_441,0,2**ADDR-1);
$readmemb("extend_file_442.mem",rom_442,0,2**ADDR-1);
$readmemb("extend_file_443.mem",rom_443,0,2**ADDR-1);
$readmemb("extend_file_444.mem",rom_444,0,2**ADDR-1);
$readmemb("extend_file_445.mem",rom_445,0,2**ADDR-1);
$readmemb("extend_file_446.mem",rom_446,0,2**ADDR-1);
$readmemb("extend_file_447.mem",rom_447,0,2**ADDR-1);
$readmemb("extend_file_448.mem",rom_448,0,2**ADDR-1);
$readmemb("extend_file_449.mem",rom_449,0,2**ADDR-1);
$readmemb("extend_file_450.mem",rom_450,0,2**ADDR-1);
$readmemb("extend_file_451.mem",rom_451,0,2**ADDR-1);
$readmemb("extend_file_452.mem",rom_452,0,2**ADDR-1);
$readmemb("extend_file_453.mem",rom_453,0,2**ADDR-1);
$readmemb("extend_file_454.mem",rom_454,0,2**ADDR-1);
$readmemb("extend_file_455.mem",rom_455,0,2**ADDR-1);
$readmemb("extend_file_456.mem",rom_456,0,2**ADDR-1);
$readmemb("extend_file_457.mem",rom_457,0,2**ADDR-1);
$readmemb("extend_file_458.mem",rom_458,0,2**ADDR-1);
$readmemb("extend_file_459.mem",rom_459,0,2**ADDR-1);
$readmemb("extend_file_460.mem",rom_460,0,2**ADDR-1);
$readmemb("extend_file_461.mem",rom_461,0,2**ADDR-1);
$readmemb("extend_file_462.mem",rom_462,0,2**ADDR-1);
$readmemb("extend_file_463.mem",rom_463,0,2**ADDR-1);
$readmemb("extend_file_464.mem",rom_464,0,2**ADDR-1);
$readmemb("extend_file_465.mem",rom_465,0,2**ADDR-1);
$readmemb("extend_file_466.mem",rom_466,0,2**ADDR-1);
$readmemb("extend_file_467.mem",rom_467,0,2**ADDR-1);
$readmemb("extend_file_468.mem",rom_468,0,2**ADDR-1);
$readmemb("extend_file_469.mem",rom_469,0,2**ADDR-1);
$readmemb("extend_file_470.mem",rom_470,0,2**ADDR-1);
$readmemb("extend_file_471.mem",rom_471,0,2**ADDR-1);
$readmemb("extend_file_472.mem",rom_472,0,2**ADDR-1);
$readmemb("extend_file_473.mem",rom_473,0,2**ADDR-1);
$readmemb("extend_file_474.mem",rom_474,0,2**ADDR-1);
$readmemb("extend_file_475.mem",rom_475,0,2**ADDR-1);
$readmemb("extend_file_476.mem",rom_476,0,2**ADDR-1);
$readmemb("extend_file_477.mem",rom_477,0,2**ADDR-1);
$readmemb("extend_file_478.mem",rom_478,0,2**ADDR-1);
$readmemb("extend_file_479.mem",rom_479,0,2**ADDR-1);
$readmemb("extend_file_480.mem",rom_480,0,2**ADDR-1);
$readmemb("extend_file_481.mem",rom_481,0,2**ADDR-1);
$readmemb("extend_file_482.mem",rom_482,0,2**ADDR-1);
$readmemb("extend_file_483.mem",rom_483,0,2**ADDR-1);
$readmemb("extend_file_484.mem",rom_484,0,2**ADDR-1);
$readmemb("extend_file_485.mem",rom_485,0,2**ADDR-1);
$readmemb("extend_file_486.mem",rom_486,0,2**ADDR-1);
$readmemb("extend_file_487.mem",rom_487,0,2**ADDR-1);
$readmemb("extend_file_488.mem",rom_488,0,2**ADDR-1);
$readmemb("extend_file_489.mem",rom_489,0,2**ADDR-1);
$readmemb("extend_file_490.mem",rom_490,0,2**ADDR-1);
$readmemb("extend_file_491.mem",rom_491,0,2**ADDR-1);
$readmemb("extend_file_492.mem",rom_492,0,2**ADDR-1);
$readmemb("extend_file_493.mem",rom_493,0,2**ADDR-1);
$readmemb("extend_file_494.mem",rom_494,0,2**ADDR-1);
$readmemb("extend_file_495.mem",rom_495,0,2**ADDR-1);
$readmemb("extend_file_496.mem",rom_496,0,2**ADDR-1);
$readmemb("extend_file_497.mem",rom_497,0,2**ADDR-1);
$readmemb("extend_file_498.mem",rom_498,0,2**ADDR-1);
$readmemb("extend_file_499.mem",rom_499,0,2**ADDR-1);
$readmemb("extend_file_500.mem",rom_500,0,2**ADDR-1);
$readmemb("extend_file_501.mem",rom_501,0,2**ADDR-1);
$readmemb("extend_file_502.mem",rom_502,0,2**ADDR-1);
$readmemb("extend_file_503.mem",rom_503,0,2**ADDR-1);
$readmemb("extend_file_504.mem",rom_504,0,2**ADDR-1);
$readmemb("extend_file_505.mem",rom_505,0,2**ADDR-1);
$readmemb("extend_file_506.mem",rom_506,0,2**ADDR-1);
$readmemb("extend_file_507.mem",rom_507,0,2**ADDR-1);
$readmemb("extend_file_508.mem",rom_508,0,2**ADDR-1);
$readmemb("extend_file_509.mem",rom_509,0,2**ADDR-1);
$readmemb("extend_file_510.mem",rom_510,0,2**ADDR-1);
$readmemb("extend_file_511.mem",rom_511,0,2**ADDR-1);
$readmemb("extend_file_512.mem",rom_512,0,2**ADDR-1);
end
assign rom_out[0] = rom_1[address] ;
assign rom_out[1] = rom_2[address] ;
assign rom_out[2] = rom_3[address] ;
assign rom_out[3] = rom_4[address] ;
assign rom_out[4] = rom_5[address] ;
assign rom_out[5] = rom_6[address] ;
assign rom_out[6] = rom_7[address] ;
assign rom_out[7] = rom_8[address] ;
assign rom_out[8] = rom_9[address] ;
assign rom_out[9] = rom_10[address] ;
assign rom_out[10] = rom_11[address] ;
assign rom_out[11] = rom_12[address] ;
assign rom_out[12] = rom_13[address] ;
assign rom_out[13] = rom_14[address] ;
assign rom_out[14] = rom_15[address] ;
assign rom_out[15] = rom_16[address] ;
assign rom_out[16] = rom_17[address] ;
assign rom_out[17] = rom_18[address] ;
assign rom_out[18] = rom_19[address] ;
assign rom_out[19] = rom_20[address] ;
assign rom_out[20] = rom_21[address] ;
assign rom_out[21] = rom_22[address] ;
assign rom_out[22] = rom_23[address] ;
assign rom_out[23] = rom_24[address] ;
assign rom_out[24] = rom_25[address] ;
assign rom_out[25] = rom_26[address] ;
assign rom_out[26] = rom_27[address] ;
assign rom_out[27] = rom_28[address] ;
assign rom_out[28] = rom_29[address] ;
assign rom_out[29] = rom_30[address] ;
assign rom_out[30] = rom_31[address] ;
assign rom_out[31] = rom_32[address] ;
assign rom_out[32] = rom_33[address] ;
assign rom_out[33] = rom_34[address] ;
assign rom_out[34] = rom_35[address] ;
assign rom_out[35] = rom_36[address] ;
assign rom_out[36] = rom_37[address] ;
assign rom_out[37] = rom_38[address] ;
assign rom_out[38] = rom_39[address] ;
assign rom_out[39] = rom_40[address] ;
assign rom_out[40] = rom_41[address] ;
assign rom_out[41] = rom_42[address] ;
assign rom_out[42] = rom_43[address] ;
assign rom_out[43] = rom_44[address] ;
assign rom_out[44] = rom_45[address] ;
assign rom_out[45] = rom_46[address] ;
assign rom_out[46] = rom_47[address] ;
assign rom_out[47] = rom_48[address] ;
assign rom_out[48] = rom_49[address] ;
assign rom_out[49] = rom_50[address] ;
assign rom_out[50] = rom_51[address] ;
assign rom_out[51] = rom_52[address] ;
assign rom_out[52] = rom_53[address] ;
assign rom_out[53] = rom_54[address] ;
assign rom_out[54] = rom_55[address] ;
assign rom_out[55] = rom_56[address] ;
assign rom_out[56] = rom_57[address] ;
assign rom_out[57] = rom_58[address] ;
assign rom_out[58] = rom_59[address] ;
assign rom_out[59] = rom_60[address] ;
assign rom_out[60] = rom_61[address] ;
assign rom_out[61] = rom_62[address] ;
assign rom_out[62] = rom_63[address] ;
assign rom_out[63] = rom_64[address] ;
assign rom_out[64] = rom_65[address] ;
assign rom_out[65] = rom_66[address] ;
assign rom_out[66] = rom_67[address] ;
assign rom_out[67] = rom_68[address] ;
assign rom_out[68] = rom_69[address] ;
assign rom_out[69] = rom_70[address] ;
assign rom_out[70] = rom_71[address] ;
assign rom_out[71] = rom_72[address] ;
assign rom_out[72] = rom_73[address] ;
assign rom_out[73] = rom_74[address] ;
assign rom_out[74] = rom_75[address] ;
assign rom_out[75] = rom_76[address] ;
assign rom_out[76] = rom_77[address] ;
assign rom_out[77] = rom_78[address] ;
assign rom_out[78] = rom_79[address] ;
assign rom_out[79] = rom_80[address] ;
assign rom_out[80] = rom_81[address] ;
assign rom_out[81] = rom_82[address] ;
assign rom_out[82] = rom_83[address] ;
assign rom_out[83] = rom_84[address] ;
assign rom_out[84] = rom_85[address] ;
assign rom_out[85] = rom_86[address] ;
assign rom_out[86] = rom_87[address] ;
assign rom_out[87] = rom_88[address] ;
assign rom_out[88] = rom_89[address] ;
assign rom_out[89] = rom_90[address] ;
assign rom_out[90] = rom_91[address] ;
assign rom_out[91] = rom_92[address] ;
assign rom_out[92] = rom_93[address] ;
assign rom_out[93] = rom_94[address] ;
assign rom_out[94] = rom_95[address] ;
assign rom_out[95] = rom_96[address] ;
assign rom_out[96] = rom_97[address] ;
assign rom_out[97] = rom_98[address] ;
assign rom_out[98] = rom_99[address] ;
assign rom_out[99] = rom_100[address] ;
assign rom_out[100] = rom_101[address] ;
assign rom_out[101] = rom_102[address] ;
assign rom_out[102] = rom_103[address] ;
assign rom_out[103] = rom_104[address] ;
assign rom_out[104] = rom_105[address] ;
assign rom_out[105] = rom_106[address] ;
assign rom_out[106] = rom_107[address] ;
assign rom_out[107] = rom_108[address] ;
assign rom_out[108] = rom_109[address] ;
assign rom_out[109] = rom_110[address] ;
assign rom_out[110] = rom_111[address] ;
assign rom_out[111] = rom_112[address] ;
assign rom_out[112] = rom_113[address] ;
assign rom_out[113] = rom_114[address] ;
assign rom_out[114] = rom_115[address] ;
assign rom_out[115] = rom_116[address] ;
assign rom_out[116] = rom_117[address] ;
assign rom_out[117] = rom_118[address] ;
assign rom_out[118] = rom_119[address] ;
assign rom_out[119] = rom_120[address] ;
assign rom_out[120] = rom_121[address] ;
assign rom_out[121] = rom_122[address] ;
assign rom_out[122] = rom_123[address] ;
assign rom_out[123] = rom_124[address] ;
assign rom_out[124] = rom_125[address] ;
assign rom_out[125] = rom_126[address] ;
assign rom_out[126] = rom_127[address] ;
assign rom_out[127] = rom_128[address] ;
assign rom_out[128] = rom_129[address] ;
assign rom_out[129] = rom_130[address] ;
assign rom_out[130] = rom_131[address] ;
assign rom_out[131] = rom_132[address] ;
assign rom_out[132] = rom_133[address] ;
assign rom_out[133] = rom_134[address] ;
assign rom_out[134] = rom_135[address] ;
assign rom_out[135] = rom_136[address] ;
assign rom_out[136] = rom_137[address] ;
assign rom_out[137] = rom_138[address] ;
assign rom_out[138] = rom_139[address] ;
assign rom_out[139] = rom_140[address] ;
assign rom_out[140] = rom_141[address] ;
assign rom_out[141] = rom_142[address] ;
assign rom_out[142] = rom_143[address] ;
assign rom_out[143] = rom_144[address] ;
assign rom_out[144] = rom_145[address] ;
assign rom_out[145] = rom_146[address] ;
assign rom_out[146] = rom_147[address] ;
assign rom_out[147] = rom_148[address] ;
assign rom_out[148] = rom_149[address] ;
assign rom_out[149] = rom_150[address] ;
assign rom_out[150] = rom_151[address] ;
assign rom_out[151] = rom_152[address] ;
assign rom_out[152] = rom_153[address] ;
assign rom_out[153] = rom_154[address] ;
assign rom_out[154] = rom_155[address] ;
assign rom_out[155] = rom_156[address] ;
assign rom_out[156] = rom_157[address] ;
assign rom_out[157] = rom_158[address] ;
assign rom_out[158] = rom_159[address] ;
assign rom_out[159] = rom_160[address] ;
assign rom_out[160] = rom_161[address] ;
assign rom_out[161] = rom_162[address] ;
assign rom_out[162] = rom_163[address] ;
assign rom_out[163] = rom_164[address] ;
assign rom_out[164] = rom_165[address] ;
assign rom_out[165] = rom_166[address] ;
assign rom_out[166] = rom_167[address] ;
assign rom_out[167] = rom_168[address] ;
assign rom_out[168] = rom_169[address] ;
assign rom_out[169] = rom_170[address] ;
assign rom_out[170] = rom_171[address] ;
assign rom_out[171] = rom_172[address] ;
assign rom_out[172] = rom_173[address] ;
assign rom_out[173] = rom_174[address] ;
assign rom_out[174] = rom_175[address] ;
assign rom_out[175] = rom_176[address] ;
assign rom_out[176] = rom_177[address] ;
assign rom_out[177] = rom_178[address] ;
assign rom_out[178] = rom_179[address] ;
assign rom_out[179] = rom_180[address] ;
assign rom_out[180] = rom_181[address] ;
assign rom_out[181] = rom_182[address] ;
assign rom_out[182] = rom_183[address] ;
assign rom_out[183] = rom_184[address] ;
assign rom_out[184] = rom_185[address] ;
assign rom_out[185] = rom_186[address] ;
assign rom_out[186] = rom_187[address] ;
assign rom_out[187] = rom_188[address] ;
assign rom_out[188] = rom_189[address] ;
assign rom_out[189] = rom_190[address] ;
assign rom_out[190] = rom_191[address] ;
assign rom_out[191] = rom_192[address] ;
assign rom_out[192] = rom_193[address] ;
assign rom_out[193] = rom_194[address] ;
assign rom_out[194] = rom_195[address] ;
assign rom_out[195] = rom_196[address] ;
assign rom_out[196] = rom_197[address] ;
assign rom_out[197] = rom_198[address] ;
assign rom_out[198] = rom_199[address] ;
assign rom_out[199] = rom_200[address] ;
assign rom_out[200] = rom_201[address] ;
assign rom_out[201] = rom_202[address] ;
assign rom_out[202] = rom_203[address] ;
assign rom_out[203] = rom_204[address] ;
assign rom_out[204] = rom_205[address] ;
assign rom_out[205] = rom_206[address] ;
assign rom_out[206] = rom_207[address] ;
assign rom_out[207] = rom_208[address] ;
assign rom_out[208] = rom_209[address] ;
assign rom_out[209] = rom_210[address] ;
assign rom_out[210] = rom_211[address] ;
assign rom_out[211] = rom_212[address] ;
assign rom_out[212] = rom_213[address] ;
assign rom_out[213] = rom_214[address] ;
assign rom_out[214] = rom_215[address] ;
assign rom_out[215] = rom_216[address] ;
assign rom_out[216] = rom_217[address] ;
assign rom_out[217] = rom_218[address] ;
assign rom_out[218] = rom_219[address] ;
assign rom_out[219] = rom_220[address] ;
assign rom_out[220] = rom_221[address] ;
assign rom_out[221] = rom_222[address] ;
assign rom_out[222] = rom_223[address] ;
assign rom_out[223] = rom_224[address] ;
assign rom_out[224] = rom_225[address] ;
assign rom_out[225] = rom_226[address] ;
assign rom_out[226] = rom_227[address] ;
assign rom_out[227] = rom_228[address] ;
assign rom_out[228] = rom_229[address] ;
assign rom_out[229] = rom_230[address] ;
assign rom_out[230] = rom_231[address] ;
assign rom_out[231] = rom_232[address] ;
assign rom_out[232] = rom_233[address] ;
assign rom_out[233] = rom_234[address] ;
assign rom_out[234] = rom_235[address] ;
assign rom_out[235] = rom_236[address] ;
assign rom_out[236] = rom_237[address] ;
assign rom_out[237] = rom_238[address] ;
assign rom_out[238] = rom_239[address] ;
assign rom_out[239] = rom_240[address] ;
assign rom_out[240] = rom_241[address] ;
assign rom_out[241] = rom_242[address] ;
assign rom_out[242] = rom_243[address] ;
assign rom_out[243] = rom_244[address] ;
assign rom_out[244] = rom_245[address] ;
assign rom_out[245] = rom_246[address] ;
assign rom_out[246] = rom_247[address] ;
assign rom_out[247] = rom_248[address] ;
assign rom_out[248] = rom_249[address] ;
assign rom_out[249] = rom_250[address] ;
assign rom_out[250] = rom_251[address] ;
assign rom_out[251] = rom_252[address] ;
assign rom_out[252] = rom_253[address] ;
assign rom_out[253] = rom_254[address] ;
assign rom_out[254] = rom_255[address] ;
assign rom_out[255] = rom_256[address] ;
assign rom_out[256] = rom_257[address] ;
assign rom_out[257] = rom_258[address] ;
assign rom_out[258] = rom_259[address] ;
assign rom_out[259] = rom_260[address] ;
assign rom_out[260] = rom_261[address] ;
assign rom_out[261] = rom_262[address] ;
assign rom_out[262] = rom_263[address] ;
assign rom_out[263] = rom_264[address] ;
assign rom_out[264] = rom_265[address] ;
assign rom_out[265] = rom_266[address] ;
assign rom_out[266] = rom_267[address] ;
assign rom_out[267] = rom_268[address] ;
assign rom_out[268] = rom_269[address] ;
assign rom_out[269] = rom_270[address] ;
assign rom_out[270] = rom_271[address] ;
assign rom_out[271] = rom_272[address] ;
assign rom_out[272] = rom_273[address] ;
assign rom_out[273] = rom_274[address] ;
assign rom_out[274] = rom_275[address] ;
assign rom_out[275] = rom_276[address] ;
assign rom_out[276] = rom_277[address] ;
assign rom_out[277] = rom_278[address] ;
assign rom_out[278] = rom_279[address] ;
assign rom_out[279] = rom_280[address] ;
assign rom_out[280] = rom_281[address] ;
assign rom_out[281] = rom_282[address] ;
assign rom_out[282] = rom_283[address] ;
assign rom_out[283] = rom_284[address] ;
assign rom_out[284] = rom_285[address] ;
assign rom_out[285] = rom_286[address] ;
assign rom_out[286] = rom_287[address] ;
assign rom_out[287] = rom_288[address] ;
assign rom_out[288] = rom_289[address] ;
assign rom_out[289] = rom_290[address] ;
assign rom_out[290] = rom_291[address] ;
assign rom_out[291] = rom_292[address] ;
assign rom_out[292] = rom_293[address] ;
assign rom_out[293] = rom_294[address] ;
assign rom_out[294] = rom_295[address] ;
assign rom_out[295] = rom_296[address] ;
assign rom_out[296] = rom_297[address] ;
assign rom_out[297] = rom_298[address] ;
assign rom_out[298] = rom_299[address] ;
assign rom_out[299] = rom_300[address] ;
assign rom_out[300] = rom_301[address] ;
assign rom_out[301] = rom_302[address] ;
assign rom_out[302] = rom_303[address] ;
assign rom_out[303] = rom_304[address] ;
assign rom_out[304] = rom_305[address] ;
assign rom_out[305] = rom_306[address] ;
assign rom_out[306] = rom_307[address] ;
assign rom_out[307] = rom_308[address] ;
assign rom_out[308] = rom_309[address] ;
assign rom_out[309] = rom_310[address] ;
assign rom_out[310] = rom_311[address] ;
assign rom_out[311] = rom_312[address] ;
assign rom_out[312] = rom_313[address] ;
assign rom_out[313] = rom_314[address] ;
assign rom_out[314] = rom_315[address] ;
assign rom_out[315] = rom_316[address] ;
assign rom_out[316] = rom_317[address] ;
assign rom_out[317] = rom_318[address] ;
assign rom_out[318] = rom_319[address] ;
assign rom_out[319] = rom_320[address] ;
assign rom_out[320] = rom_321[address] ;
assign rom_out[321] = rom_322[address] ;
assign rom_out[322] = rom_323[address] ;
assign rom_out[323] = rom_324[address] ;
assign rom_out[324] = rom_325[address] ;
assign rom_out[325] = rom_326[address] ;
assign rom_out[326] = rom_327[address] ;
assign rom_out[327] = rom_328[address] ;
assign rom_out[328] = rom_329[address] ;
assign rom_out[329] = rom_330[address] ;
assign rom_out[330] = rom_331[address] ;
assign rom_out[331] = rom_332[address] ;
assign rom_out[332] = rom_333[address] ;
assign rom_out[333] = rom_334[address] ;
assign rom_out[334] = rom_335[address] ;
assign rom_out[335] = rom_336[address] ;
assign rom_out[336] = rom_337[address] ;
assign rom_out[337] = rom_338[address] ;
assign rom_out[338] = rom_339[address] ;
assign rom_out[339] = rom_340[address] ;
assign rom_out[340] = rom_341[address] ;
assign rom_out[341] = rom_342[address] ;
assign rom_out[342] = rom_343[address] ;
assign rom_out[343] = rom_344[address] ;
assign rom_out[344] = rom_345[address] ;
assign rom_out[345] = rom_346[address] ;
assign rom_out[346] = rom_347[address] ;
assign rom_out[347] = rom_348[address] ;
assign rom_out[348] = rom_349[address] ;
assign rom_out[349] = rom_350[address] ;
assign rom_out[350] = rom_351[address] ;
assign rom_out[351] = rom_352[address] ;
assign rom_out[352] = rom_353[address] ;
assign rom_out[353] = rom_354[address] ;
assign rom_out[354] = rom_355[address] ;
assign rom_out[355] = rom_356[address] ;
assign rom_out[356] = rom_357[address] ;
assign rom_out[357] = rom_358[address] ;
assign rom_out[358] = rom_359[address] ;
assign rom_out[359] = rom_360[address] ;
assign rom_out[360] = rom_361[address] ;
assign rom_out[361] = rom_362[address] ;
assign rom_out[362] = rom_363[address] ;
assign rom_out[363] = rom_364[address] ;
assign rom_out[364] = rom_365[address] ;
assign rom_out[365] = rom_366[address] ;
assign rom_out[366] = rom_367[address] ;
assign rom_out[367] = rom_368[address] ;
assign rom_out[368] = rom_369[address] ;
assign rom_out[369] = rom_370[address] ;
assign rom_out[370] = rom_371[address] ;
assign rom_out[371] = rom_372[address] ;
assign rom_out[372] = rom_373[address] ;
assign rom_out[373] = rom_374[address] ;
assign rom_out[374] = rom_375[address] ;
assign rom_out[375] = rom_376[address] ;
assign rom_out[376] = rom_377[address] ;
assign rom_out[377] = rom_378[address] ;
assign rom_out[378] = rom_379[address] ;
assign rom_out[379] = rom_380[address] ;
assign rom_out[380] = rom_381[address] ;
assign rom_out[381] = rom_382[address] ;
assign rom_out[382] = rom_383[address] ;
assign rom_out[383] = rom_384[address] ;
assign rom_out[384] = rom_385[address] ;
assign rom_out[385] = rom_386[address] ;
assign rom_out[386] = rom_387[address] ;
assign rom_out[387] = rom_388[address] ;
assign rom_out[388] = rom_389[address] ;
assign rom_out[389] = rom_390[address] ;
assign rom_out[390] = rom_391[address] ;
assign rom_out[391] = rom_392[address] ;
assign rom_out[392] = rom_393[address] ;
assign rom_out[393] = rom_394[address] ;
assign rom_out[394] = rom_395[address] ;
assign rom_out[395] = rom_396[address] ;
assign rom_out[396] = rom_397[address] ;
assign rom_out[397] = rom_398[address] ;
assign rom_out[398] = rom_399[address] ;
assign rom_out[399] = rom_400[address] ;
assign rom_out[400] = rom_401[address] ;
assign rom_out[401] = rom_402[address] ;
assign rom_out[402] = rom_403[address] ;
assign rom_out[403] = rom_404[address] ;
assign rom_out[404] = rom_405[address] ;
assign rom_out[405] = rom_406[address] ;
assign rom_out[406] = rom_407[address] ;
assign rom_out[407] = rom_408[address] ;
assign rom_out[408] = rom_409[address] ;
assign rom_out[409] = rom_410[address] ;
assign rom_out[410] = rom_411[address] ;
assign rom_out[411] = rom_412[address] ;
assign rom_out[412] = rom_413[address] ;
assign rom_out[413] = rom_414[address] ;
assign rom_out[414] = rom_415[address] ;
assign rom_out[415] = rom_416[address] ;
assign rom_out[416] = rom_417[address] ;
assign rom_out[417] = rom_418[address] ;
assign rom_out[418] = rom_419[address] ;
assign rom_out[419] = rom_420[address] ;
assign rom_out[420] = rom_421[address] ;
assign rom_out[421] = rom_422[address] ;
assign rom_out[422] = rom_423[address] ;
assign rom_out[423] = rom_424[address] ;
assign rom_out[424] = rom_425[address] ;
assign rom_out[425] = rom_426[address] ;
assign rom_out[426] = rom_427[address] ;
assign rom_out[427] = rom_428[address] ;
assign rom_out[428] = rom_429[address] ;
assign rom_out[429] = rom_430[address] ;
assign rom_out[430] = rom_431[address] ;
assign rom_out[431] = rom_432[address] ;
assign rom_out[432] = rom_433[address] ;
assign rom_out[433] = rom_434[address] ;
assign rom_out[434] = rom_435[address] ;
assign rom_out[435] = rom_436[address] ;
assign rom_out[436] = rom_437[address] ;
assign rom_out[437] = rom_438[address] ;
assign rom_out[438] = rom_439[address] ;
assign rom_out[439] = rom_440[address] ;
assign rom_out[440] = rom_441[address] ;
assign rom_out[441] = rom_442[address] ;
assign rom_out[442] = rom_443[address] ;
assign rom_out[443] = rom_444[address] ;
assign rom_out[444] = rom_445[address] ;
assign rom_out[445] = rom_446[address] ;
assign rom_out[446] = rom_447[address] ;
assign rom_out[447] = rom_448[address] ;
assign rom_out[448] = rom_449[address] ;
assign rom_out[449] = rom_450[address] ;
assign rom_out[450] = rom_451[address] ;
assign rom_out[451] = rom_452[address] ;
assign rom_out[452] = rom_453[address] ;
assign rom_out[453] = rom_454[address] ;
assign rom_out[454] = rom_455[address] ;
assign rom_out[455] = rom_456[address] ;
assign rom_out[456] = rom_457[address] ;
assign rom_out[457] = rom_458[address] ;
assign rom_out[458] = rom_459[address] ;
assign rom_out[459] = rom_460[address] ;
assign rom_out[460] = rom_461[address] ;
assign rom_out[461] = rom_462[address] ;
assign rom_out[462] = rom_463[address] ;
assign rom_out[463] = rom_464[address] ;
assign rom_out[464] = rom_465[address] ;
assign rom_out[465] = rom_466[address] ;
assign rom_out[466] = rom_467[address] ;
assign rom_out[467] = rom_468[address] ;
assign rom_out[468] = rom_469[address] ;
assign rom_out[469] = rom_470[address] ;
assign rom_out[470] = rom_471[address] ;
assign rom_out[471] = rom_472[address] ;
assign rom_out[472] = rom_473[address] ;
assign rom_out[473] = rom_474[address] ;
assign rom_out[474] = rom_475[address] ;
assign rom_out[475] = rom_476[address] ;
assign rom_out[476] = rom_477[address] ;
assign rom_out[477] = rom_478[address] ;
assign rom_out[478] = rom_479[address] ;
assign rom_out[479] = rom_480[address] ;
assign rom_out[480] = rom_481[address] ;
assign rom_out[481] = rom_482[address] ;
assign rom_out[482] = rom_483[address] ;
assign rom_out[483] = rom_484[address] ;
assign rom_out[484] = rom_485[address] ;
assign rom_out[485] = rom_486[address] ;
assign rom_out[486] = rom_487[address] ;
assign rom_out[487] = rom_488[address] ;
assign rom_out[488] = rom_489[address] ;
assign rom_out[489] = rom_490[address] ;
assign rom_out[490] = rom_491[address] ;
assign rom_out[491] = rom_492[address] ;
assign rom_out[492] = rom_493[address] ;
assign rom_out[493] = rom_494[address] ;
assign rom_out[494] = rom_495[address] ;
assign rom_out[495] = rom_496[address] ;
assign rom_out[496] = rom_497[address] ;
assign rom_out[497] = rom_498[address] ;
assign rom_out[498] = rom_499[address] ;
assign rom_out[499] = rom_500[address] ;
assign rom_out[500] = rom_501[address] ;
assign rom_out[501] = rom_502[address] ;
assign rom_out[502] = rom_503[address] ;
assign rom_out[503] = rom_504[address] ;
assign rom_out[504] = rom_505[address] ;
assign rom_out[505] = rom_506[address] ;
assign rom_out[506] = rom_507[address] ;
assign rom_out[507] = rom_508[address] ;
assign rom_out[508] = rom_509[address] ;
assign rom_out[509] = rom_510[address] ;
assign rom_out[510] = rom_511[address] ;
assign rom_out[511] = rom_512[address] ;
endmodule
