
module biasing_rom (
	output [15:0] bias_mem [0:112-1]
);

reg [16-1:0] bias_reg_0 = 16'b0000000011001111;
reg [16-1:0] bias_reg_1 = 16'b1000000100101111;
reg [16-1:0] bias_reg_2 = 16'b0000000010100101;
reg [16-1:0] bias_reg_3 = 16'b0000000001110111;
reg [16-1:0] bias_reg_4 = 16'b1000000111100000;
reg [16-1:0] bias_reg_5 = 16'b1000000010100100;
reg [16-1:0] bias_reg_6 = 16'b0000000011111111;
reg [16-1:0] bias_reg_7 = 16'b1000001011000011;
reg [16-1:0] bias_reg_8 = 16'b1000000100000101;
reg [16-1:0] bias_reg_9 = 16'b1000000000111000;
reg [16-1:0] bias_reg_10 = 16'b0000000001110000;
reg [16-1:0] bias_reg_11 = 16'b1000000010010100;
reg [16-1:0] bias_reg_12 = 16'b1000000001001111;
reg [16-1:0] bias_reg_13 = 16'b0000000010010101;
reg [16-1:0] bias_reg_14 = 16'b1000000010011101;
reg [16-1:0] bias_reg_15 = 16'b1000000001001000;
reg [16-1:0] bias_reg_16 = 16'b0000000001111000;
reg [16-1:0] bias_reg_17 = 16'b1000000010100000;
reg [16-1:0] bias_reg_18 = 16'b0000000010000001;
reg [16-1:0] bias_reg_19 = 16'b0000000010100000;
reg [16-1:0] bias_reg_20 = 16'b0000000100010110;
reg [16-1:0] bias_reg_21 = 16'b1000011000011000;
reg [16-1:0] bias_reg_22 = 16'b1000000011010011;
reg [16-1:0] bias_reg_23 = 16'b0000000001111011;
reg [16-1:0] bias_reg_24 = 16'b0000000101010010;
reg [16-1:0] bias_reg_25 = 16'b0000000100001010;
reg [16-1:0] bias_reg_26 = 16'b1000000001100100;
reg [16-1:0] bias_reg_27 = 16'b0000000000010001;
reg [16-1:0] bias_reg_28 = 16'b0000000000010010;
reg [16-1:0] bias_reg_29 = 16'b0000000010011001;
reg [16-1:0] bias_reg_30 = 16'b1000000010110000;
reg [16-1:0] bias_reg_31 = 16'b0000000001000010;
reg [16-1:0] bias_reg_32 = 16'b1000000001011000;
reg [16-1:0] bias_reg_33 = 16'b0000000000110000;
reg [16-1:0] bias_reg_34 = 16'b1000000101010000;
reg [16-1:0] bias_reg_35 = 16'b1000000110001010;
reg [16-1:0] bias_reg_36 = 16'b1000000011110111;
reg [16-1:0] bias_reg_37 = 16'b1000101111111101;
reg [16-1:0] bias_reg_38 = 16'b1000001001010111;
reg [16-1:0] bias_reg_39 = 16'b0000000000000001;
reg [16-1:0] bias_reg_40 = 16'b1000000110011010;
reg [16-1:0] bias_reg_41 = 16'b0000000010100010;
reg [16-1:0] bias_reg_42 = 16'b0000000101010101;
reg [16-1:0] bias_reg_43 = 16'b1000000110000010;
reg [16-1:0] bias_reg_44 = 16'b0000000110111010;
reg [16-1:0] bias_reg_45 = 16'b0000000001101111;
reg [16-1:0] bias_reg_46 = 16'b0000000000110000;
reg [16-1:0] bias_reg_47 = 16'b1000000000010111;
reg [16-1:0] bias_reg_48 = 16'b1000000010100011;
reg [16-1:0] bias_reg_49 = 16'b1000000000001110;
reg [16-1:0] bias_reg_50 = 16'b1000000101000010;
reg [16-1:0] bias_reg_51 = 16'b1000000111110101;
reg [16-1:0] bias_reg_52 = 16'b1000000001111111;
reg [16-1:0] bias_reg_53 = 16'b0000000000000101;
reg [16-1:0] bias_reg_54 = 16'b1000000000111100;
reg [16-1:0] bias_reg_55 = 16'b0000000001100001;
reg [16-1:0] bias_reg_56 = 16'b0000000000111011;
reg [16-1:0] bias_reg_57 = 16'b1000000110000011;
reg [16-1:0] bias_reg_58 = 16'b0000100100011001;
reg [16-1:0] bias_reg_59 = 16'b0000000001110101;
reg [16-1:0] bias_reg_60 = 16'b0000000000110111;
reg [16-1:0] bias_reg_61 = 16'b1000000000011110;
reg [16-1:0] bias_reg_62 = 16'b0000000001101110;
reg [16-1:0] bias_reg_63 = 16'b0000000010010001;
reg [16-1:0] bias_reg_64 = 16'b0000000100001010;
reg [16-1:0] bias_reg_65 = 16'b0000000000000100;
reg [16-1:0] bias_reg_66 = 16'b0000000001100010;
reg [16-1:0] bias_reg_67 = 16'b0000000001000000;
reg [16-1:0] bias_reg_68 = 16'b0000000011011111;
reg [16-1:0] bias_reg_69 = 16'b1000001000111110;
reg [16-1:0] bias_reg_70 = 16'b0000000000100111;
reg [16-1:0] bias_reg_71 = 16'b1000001101101001;
reg [16-1:0] bias_reg_72 = 16'b0000000100100110;
reg [16-1:0] bias_reg_73 = 16'b1000000000011011;
reg [16-1:0] bias_reg_74 = 16'b1000000000100011;
reg [16-1:0] bias_reg_75 = 16'b1000001010100010;
reg [16-1:0] bias_reg_76 = 16'b1000000001110111;
reg [16-1:0] bias_reg_77 = 16'b0000000101000110;
reg [16-1:0] bias_reg_78 = 16'b1000000011010100;
reg [16-1:0] bias_reg_79 = 16'b0000000010000011;
reg [16-1:0] bias_reg_80 = 16'b0000000010100100;
reg [16-1:0] bias_reg_81 = 16'b1000000000000101;
reg [16-1:0] bias_reg_82 = 16'b1000000010000100;
reg [16-1:0] bias_reg_83 = 16'b0000000001010111;
reg [16-1:0] bias_reg_84 = 16'b1000000000011000;
reg [16-1:0] bias_reg_85 = 16'b0000000001000000;
reg [16-1:0] bias_reg_86 = 16'b1000001011110111;
reg [16-1:0] bias_reg_87 = 16'b1000000100000000;
reg [16-1:0] bias_reg_88 = 16'b0000000100010001;
reg [16-1:0] bias_reg_89 = 16'b0000000001100011;
reg [16-1:0] bias_reg_90 = 16'b0000000000010010;
reg [16-1:0] bias_reg_91 = 16'b0000000010000011;
reg [16-1:0] bias_reg_92 = 16'b0000000011101010;
reg [16-1:0] bias_reg_93 = 16'b1000000110000010;
reg [16-1:0] bias_reg_94 = 16'b1000000100001010;
reg [16-1:0] bias_reg_95 = 16'b1000000010010111;
reg [16-1:0] bias_reg_96 = 16'b1000000001011110;
reg [16-1:0] bias_reg_97 = 16'b1000000000010010;
reg [16-1:0] bias_reg_98 = 16'b1000001010011100;
reg [16-1:0] bias_reg_99 = 16'b0000000011011100;
reg [16-1:0] bias_reg_100 = 16'b1000000001010101;
reg [16-1:0] bias_reg_101 = 16'b0000000011001111;
reg [16-1:0] bias_reg_102 = 16'b0000000010010110;
reg [16-1:0] bias_reg_103 = 16'b0000000101000000;
reg [16-1:0] bias_reg_104 = 16'b0000000001101110;
reg [16-1:0] bias_reg_105 = 16'b1000001000001010;
reg [16-1:0] bias_reg_106 = 16'b0000000011110001;
reg [16-1:0] bias_reg_107 = 16'b1000001100000011;
reg [16-1:0] bias_reg_108 = 16'b1000000001100110;
reg [16-1:0] bias_reg_109 = 16'b0000000001111001;
reg [16-1:0] bias_reg_110 = 16'b1000000000101100;
reg [16-1:0] bias_reg_111 = 16'b1000000010100000;
assign bias_mem[0] = bias_reg_0;
assign bias_mem[1] = bias_reg_1;
assign bias_mem[2] = bias_reg_2;
assign bias_mem[3] = bias_reg_3;
assign bias_mem[4] = bias_reg_4;
assign bias_mem[5] = bias_reg_5;
assign bias_mem[6] = bias_reg_6;
assign bias_mem[7] = bias_reg_7;
assign bias_mem[8] = bias_reg_8;
assign bias_mem[9] = bias_reg_9;
assign bias_mem[10] = bias_reg_10;
assign bias_mem[11] = bias_reg_11;
assign bias_mem[12] = bias_reg_12;
assign bias_mem[13] = bias_reg_13;
assign bias_mem[14] = bias_reg_14;
assign bias_mem[15] = bias_reg_15;
assign bias_mem[16] = bias_reg_16;
assign bias_mem[17] = bias_reg_17;
assign bias_mem[18] = bias_reg_18;
assign bias_mem[19] = bias_reg_19;
assign bias_mem[20] = bias_reg_20;
assign bias_mem[21] = bias_reg_21;
assign bias_mem[22] = bias_reg_22;
assign bias_mem[23] = bias_reg_23;
assign bias_mem[24] = bias_reg_24;
assign bias_mem[25] = bias_reg_25;
assign bias_mem[26] = bias_reg_26;
assign bias_mem[27] = bias_reg_27;
assign bias_mem[28] = bias_reg_28;
assign bias_mem[29] = bias_reg_29;
assign bias_mem[30] = bias_reg_30;
assign bias_mem[31] = bias_reg_31;
assign bias_mem[32] = bias_reg_32;
assign bias_mem[33] = bias_reg_33;
assign bias_mem[34] = bias_reg_34;
assign bias_mem[35] = bias_reg_35;
assign bias_mem[36] = bias_reg_36;
assign bias_mem[37] = bias_reg_37;
assign bias_mem[38] = bias_reg_38;
assign bias_mem[39] = bias_reg_39;
assign bias_mem[40] = bias_reg_40;
assign bias_mem[41] = bias_reg_41;
assign bias_mem[42] = bias_reg_42;
assign bias_mem[43] = bias_reg_43;
assign bias_mem[44] = bias_reg_44;
assign bias_mem[45] = bias_reg_45;
assign bias_mem[46] = bias_reg_46;
assign bias_mem[47] = bias_reg_47;
assign bias_mem[48] = bias_reg_48;
assign bias_mem[49] = bias_reg_49;
assign bias_mem[50] = bias_reg_50;
assign bias_mem[51] = bias_reg_51;
assign bias_mem[52] = bias_reg_52;
assign bias_mem[53] = bias_reg_53;
assign bias_mem[54] = bias_reg_54;
assign bias_mem[55] = bias_reg_55;
assign bias_mem[56] = bias_reg_56;
assign bias_mem[57] = bias_reg_57;
assign bias_mem[58] = bias_reg_58;
assign bias_mem[59] = bias_reg_59;
assign bias_mem[60] = bias_reg_60;
assign bias_mem[61] = bias_reg_61;
assign bias_mem[62] = bias_reg_62;
assign bias_mem[63] = bias_reg_63;
assign bias_mem[64] = bias_reg_64;
assign bias_mem[65] = bias_reg_65;
assign bias_mem[66] = bias_reg_66;
assign bias_mem[67] = bias_reg_67;
assign bias_mem[68] = bias_reg_68;
assign bias_mem[69] = bias_reg_69;
assign bias_mem[70] = bias_reg_70;
assign bias_mem[71] = bias_reg_71;
assign bias_mem[72] = bias_reg_72;
assign bias_mem[73] = bias_reg_73;
assign bias_mem[74] = bias_reg_74;
assign bias_mem[75] = bias_reg_75;
assign bias_mem[76] = bias_reg_76;
assign bias_mem[77] = bias_reg_77;
assign bias_mem[78] = bias_reg_78;
assign bias_mem[79] = bias_reg_79;
assign bias_mem[80] = bias_reg_80;
assign bias_mem[81] = bias_reg_81;
assign bias_mem[82] = bias_reg_82;
assign bias_mem[83] = bias_reg_83;
assign bias_mem[84] = bias_reg_84;
assign bias_mem[85] = bias_reg_85;
assign bias_mem[86] = bias_reg_86;
assign bias_mem[87] = bias_reg_87;
assign bias_mem[88] = bias_reg_88;
assign bias_mem[89] = bias_reg_89;
assign bias_mem[90] = bias_reg_90;
assign bias_mem[91] = bias_reg_91;
assign bias_mem[92] = bias_reg_92;
assign bias_mem[93] = bias_reg_93;
assign bias_mem[94] = bias_reg_94;
assign bias_mem[95] = bias_reg_95;
assign bias_mem[96] = bias_reg_96;
assign bias_mem[97] = bias_reg_97;
assign bias_mem[98] = bias_reg_98;
assign bias_mem[99] = bias_reg_99;
assign bias_mem[100] = bias_reg_100;
assign bias_mem[101] = bias_reg_101;
assign bias_mem[102] = bias_reg_102;
assign bias_mem[103] = bias_reg_103;
assign bias_mem[104] = bias_reg_104;
assign bias_mem[105] = bias_reg_105;
assign bias_mem[106] = bias_reg_106;
assign bias_mem[107] = bias_reg_107;
assign bias_mem[108] = bias_reg_108;
assign bias_mem[109] = bias_reg_109;
assign bias_mem[110] = bias_reg_110;
assign bias_mem[111] = bias_reg_111;
endmodule
