
module biasing_rom (
	output [15:0] bias_mem [0:64-1]
);

reg [16-1:0] bias_reg_0 = 16'b1000000000000001;
reg [16-1:0] bias_reg_1 = 16'b1000000000101110;
reg [16-1:0] bias_reg_2 = 16'b0000000000101000;
reg [16-1:0] bias_reg_3 = 16'b0000000011101111;
reg [16-1:0] bias_reg_4 = 16'b1000000001001111;
reg [16-1:0] bias_reg_5 = 16'b1000000001000010;
reg [16-1:0] bias_reg_6 = 16'b1000000000100011;
reg [16-1:0] bias_reg_7 = 16'b0000000000001100;
reg [16-1:0] bias_reg_8 = 16'b1000000000001101;
reg [16-1:0] bias_reg_9 = 16'b0000000000000000;
reg [16-1:0] bias_reg_10 = 16'b1000000000111011;
reg [16-1:0] bias_reg_11 = 16'b1000000001010100;
reg [16-1:0] bias_reg_12 = 16'b1000000001000100;
reg [16-1:0] bias_reg_13 = 16'b0000000000001011;
reg [16-1:0] bias_reg_14 = 16'b0000000001110110;
reg [16-1:0] bias_reg_15 = 16'b1000000000110111;
reg [16-1:0] bias_reg_16 = 16'b1000000000100000;
reg [16-1:0] bias_reg_17 = 16'b1000000001001110;
reg [16-1:0] bias_reg_18 = 16'b1000000000011000;
reg [16-1:0] bias_reg_19 = 16'b1000000000000001;
reg [16-1:0] bias_reg_20 = 16'b0000000011000010;
reg [16-1:0] bias_reg_21 = 16'b0000000100001101;
reg [16-1:0] bias_reg_22 = 16'b1000000010001010;
reg [16-1:0] bias_reg_23 = 16'b0000000001010101;
reg [16-1:0] bias_reg_24 = 16'b1000000001000011;
reg [16-1:0] bias_reg_25 = 16'b1000000010100010;
reg [16-1:0] bias_reg_26 = 16'b0000000000010100;
reg [16-1:0] bias_reg_27 = 16'b1000000001011010;
reg [16-1:0] bias_reg_28 = 16'b1000000000100101;
reg [16-1:0] bias_reg_29 = 16'b1000000001101100;
reg [16-1:0] bias_reg_30 = 16'b1000000000000001;
reg [16-1:0] bias_reg_31 = 16'b0000000000000000;
reg [16-1:0] bias_reg_32 = 16'b0000000011110000;
reg [16-1:0] bias_reg_33 = 16'b1000000011001101;
reg [16-1:0] bias_reg_34 = 16'b1000000001000011;
reg [16-1:0] bias_reg_35 = 16'b0000000000000000;
reg [16-1:0] bias_reg_36 = 16'b0000000000000000;
reg [16-1:0] bias_reg_37 = 16'b1000000011000100;
reg [16-1:0] bias_reg_38 = 16'b0000000000110111;
reg [16-1:0] bias_reg_39 = 16'b1000000000000001;
reg [16-1:0] bias_reg_40 = 16'b1000000001111000;
reg [16-1:0] bias_reg_41 = 16'b1000000001110010;
reg [16-1:0] bias_reg_42 = 16'b0000000001000001;
reg [16-1:0] bias_reg_43 = 16'b1000000000111110;
reg [16-1:0] bias_reg_44 = 16'b0000000010101101;
reg [16-1:0] bias_reg_45 = 16'b1000000010011010;
reg [16-1:0] bias_reg_46 = 16'b1000000001100111;
reg [16-1:0] bias_reg_47 = 16'b1000000000000001;
reg [16-1:0] bias_reg_48 = 16'b1000000000000001;
reg [16-1:0] bias_reg_49 = 16'b1000000000111000;
reg [16-1:0] bias_reg_50 = 16'b1000000001000100;
reg [16-1:0] bias_reg_51 = 16'b1000000001000000;
reg [16-1:0] bias_reg_52 = 16'b1000000001101111;
reg [16-1:0] bias_reg_53 = 16'b1000000000000001;
reg [16-1:0] bias_reg_54 = 16'b0000000001111011;
reg [16-1:0] bias_reg_55 = 16'b1000000000000001;
reg [16-1:0] bias_reg_56 = 16'b0000000000000000;
reg [16-1:0] bias_reg_57 = 16'b1000000001011110;
reg [16-1:0] bias_reg_58 = 16'b0000000010000101;
reg [16-1:0] bias_reg_59 = 16'b1000000000001010;
reg [16-1:0] bias_reg_60 = 16'b1000000001011000;
reg [16-1:0] bias_reg_61 = 16'b1000000000110000;
reg [16-1:0] bias_reg_62 = 16'b1000000001000111;
reg [16-1:0] bias_reg_63 = 16'b1000000000000001;
assign bias_mem[0] = bias_reg_0;
assign bias_mem[1] = bias_reg_1;
assign bias_mem[2] = bias_reg_2;
assign bias_mem[3] = bias_reg_3;
assign bias_mem[4] = bias_reg_4;
assign bias_mem[5] = bias_reg_5;
assign bias_mem[6] = bias_reg_6;
assign bias_mem[7] = bias_reg_7;
assign bias_mem[8] = bias_reg_8;
assign bias_mem[9] = bias_reg_9;
assign bias_mem[10] = bias_reg_10;
assign bias_mem[11] = bias_reg_11;
assign bias_mem[12] = bias_reg_12;
assign bias_mem[13] = bias_reg_13;
assign bias_mem[14] = bias_reg_14;
assign bias_mem[15] = bias_reg_15;
assign bias_mem[16] = bias_reg_16;
assign bias_mem[17] = bias_reg_17;
assign bias_mem[18] = bias_reg_18;
assign bias_mem[19] = bias_reg_19;
assign bias_mem[20] = bias_reg_20;
assign bias_mem[21] = bias_reg_21;
assign bias_mem[22] = bias_reg_22;
assign bias_mem[23] = bias_reg_23;
assign bias_mem[24] = bias_reg_24;
assign bias_mem[25] = bias_reg_25;
assign bias_mem[26] = bias_reg_26;
assign bias_mem[27] = bias_reg_27;
assign bias_mem[28] = bias_reg_28;
assign bias_mem[29] = bias_reg_29;
assign bias_mem[30] = bias_reg_30;
assign bias_mem[31] = bias_reg_31;
assign bias_mem[32] = bias_reg_32;
assign bias_mem[33] = bias_reg_33;
assign bias_mem[34] = bias_reg_34;
assign bias_mem[35] = bias_reg_35;
assign bias_mem[36] = bias_reg_36;
assign bias_mem[37] = bias_reg_37;
assign bias_mem[38] = bias_reg_38;
assign bias_mem[39] = bias_reg_39;
assign bias_mem[40] = bias_reg_40;
assign bias_mem[41] = bias_reg_41;
assign bias_mem[42] = bias_reg_42;
assign bias_mem[43] = bias_reg_43;
assign bias_mem[44] = bias_reg_44;
assign bias_mem[45] = bias_reg_45;
assign bias_mem[46] = bias_reg_46;
assign bias_mem[47] = bias_reg_47;
assign bias_mem[48] = bias_reg_48;
assign bias_mem[49] = bias_reg_49;
assign bias_mem[50] = bias_reg_50;
assign bias_mem[51] = bias_reg_51;
assign bias_mem[52] = bias_reg_52;
assign bias_mem[53] = bias_reg_53;
assign bias_mem[54] = bias_reg_54;
assign bias_mem[55] = bias_reg_55;
assign bias_mem[56] = bias_reg_56;
assign bias_mem[57] = bias_reg_57;
assign bias_mem[58] = bias_reg_58;
assign bias_mem[59] = bias_reg_59;
assign bias_mem[60] = bias_reg_60;
assign bias_mem[61] = bias_reg_61;
assign bias_mem[62] = bias_reg_62;
assign bias_mem[63] = bias_reg_63;
endmodule
