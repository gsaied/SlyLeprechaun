
module biasing_rom (
	output [15:0] bias_mem [0:32-1]
);

reg [16-1:0] bias_reg_0 = 16'b1000000000101110;
reg [16-1:0] bias_reg_1 = 16'b0000000001001000;
reg [16-1:0] bias_reg_2 = 16'b0000000001010010;
reg [16-1:0] bias_reg_3 = 16'b1000000010010110;
reg [16-1:0] bias_reg_4 = 16'b0000000000011000;
reg [16-1:0] bias_reg_5 = 16'b0000000001100101;
reg [16-1:0] bias_reg_6 = 16'b0000000010011010;
reg [16-1:0] bias_reg_7 = 16'b1000000000000111;
reg [16-1:0] bias_reg_8 = 16'b1000000010000011;
reg [16-1:0] bias_reg_9 = 16'b0000000000000111;
reg [16-1:0] bias_reg_10 = 16'b0000000000011101;
reg [16-1:0] bias_reg_11 = 16'b1000000001001010;
reg [16-1:0] bias_reg_12 = 16'b1000001010100001;
reg [16-1:0] bias_reg_13 = 16'b0000001010000000;
reg [16-1:0] bias_reg_14 = 16'b1000000000011010;
reg [16-1:0] bias_reg_15 = 16'b0000000110111001;
reg [16-1:0] bias_reg_16 = 16'b0000000010011110;
reg [16-1:0] bias_reg_17 = 16'b1000000001101101;
reg [16-1:0] bias_reg_18 = 16'b0000000000010011;
reg [16-1:0] bias_reg_19 = 16'b0000000001010011;
reg [16-1:0] bias_reg_20 = 16'b0000000000011101;
reg [16-1:0] bias_reg_21 = 16'b0000000001000010;
reg [16-1:0] bias_reg_22 = 16'b0000000001011010;
reg [16-1:0] bias_reg_23 = 16'b0000000000001000;
reg [16-1:0] bias_reg_24 = 16'b0000000000001101;
reg [16-1:0] bias_reg_25 = 16'b1000000001000011;
reg [16-1:0] bias_reg_26 = 16'b0000000011010100;
reg [16-1:0] bias_reg_27 = 16'b0000000000000111;
reg [16-1:0] bias_reg_28 = 16'b0000000000110111;
reg [16-1:0] bias_reg_29 = 16'b1000000000110101;
reg [16-1:0] bias_reg_30 = 16'b0000000000101010;
reg [16-1:0] bias_reg_31 = 16'b1000000000000110;
assign bias_mem[0] = bias_reg_0;
assign bias_mem[1] = bias_reg_1;
assign bias_mem[2] = bias_reg_2;
assign bias_mem[3] = bias_reg_3;
assign bias_mem[4] = bias_reg_4;
assign bias_mem[5] = bias_reg_5;
assign bias_mem[6] = bias_reg_6;
assign bias_mem[7] = bias_reg_7;
assign bias_mem[8] = bias_reg_8;
assign bias_mem[9] = bias_reg_9;
assign bias_mem[10] = bias_reg_10;
assign bias_mem[11] = bias_reg_11;
assign bias_mem[12] = bias_reg_12;
assign bias_mem[13] = bias_reg_13;
assign bias_mem[14] = bias_reg_14;
assign bias_mem[15] = bias_reg_15;
assign bias_mem[16] = bias_reg_16;
assign bias_mem[17] = bias_reg_17;
assign bias_mem[18] = bias_reg_18;
assign bias_mem[19] = bias_reg_19;
assign bias_mem[20] = bias_reg_20;
assign bias_mem[21] = bias_reg_21;
assign bias_mem[22] = bias_reg_22;
assign bias_mem[23] = bias_reg_23;
assign bias_mem[24] = bias_reg_24;
assign bias_mem[25] = bias_reg_25;
assign bias_mem[26] = bias_reg_26;
assign bias_mem[27] = bias_reg_27;
assign bias_mem[28] = bias_reg_28;
assign bias_mem[29] = bias_reg_29;
assign bias_mem[30] = bias_reg_30;
assign bias_mem[31] = bias_reg_31;
endmodule
