
module biasing_rom (
	output [15:0] bias_mem [0:368-1]
);

reg [16-1:0] bias_reg_0 = 16'b0000000000101101;
reg [16-1:0] bias_reg_1 = 16'b0000000010011011;
reg [16-1:0] bias_reg_2 = 16'b0000000001011100;
reg [16-1:0] bias_reg_3 = 16'b0000000001100101;
reg [16-1:0] bias_reg_4 = 16'b0000000010100101;
reg [16-1:0] bias_reg_5 = 16'b0000000001000010;
reg [16-1:0] bias_reg_6 = 16'b0000000010010000;
reg [16-1:0] bias_reg_7 = 16'b0000000000110011;
reg [16-1:0] bias_reg_8 = 16'b0000000001011000;
reg [16-1:0] bias_reg_9 = 16'b0000000001001111;
reg [16-1:0] bias_reg_10 = 16'b0000000001010111;
reg [16-1:0] bias_reg_11 = 16'b0000000001001111;
reg [16-1:0] bias_reg_12 = 16'b0000000010100010;
reg [16-1:0] bias_reg_13 = 16'b0000000001100100;
reg [16-1:0] bias_reg_14 = 16'b0000000000101100;
reg [16-1:0] bias_reg_15 = 16'b0000000000111001;
reg [16-1:0] bias_reg_16 = 16'b0000000000101000;
reg [16-1:0] bias_reg_17 = 16'b0000000001011001;
reg [16-1:0] bias_reg_18 = 16'b0000000011001001;
reg [16-1:0] bias_reg_19 = 16'b0000000000101110;
reg [16-1:0] bias_reg_20 = 16'b0000000001101101;
reg [16-1:0] bias_reg_21 = 16'b0000000100001100;
reg [16-1:0] bias_reg_22 = 16'b0000000001000011;
reg [16-1:0] bias_reg_23 = 16'b0000000010001110;
reg [16-1:0] bias_reg_24 = 16'b0000000010000010;
reg [16-1:0] bias_reg_25 = 16'b0000000001001000;
reg [16-1:0] bias_reg_26 = 16'b0000000001001000;
reg [16-1:0] bias_reg_27 = 16'b0000000001001101;
reg [16-1:0] bias_reg_28 = 16'b0000000001010000;
reg [16-1:0] bias_reg_29 = 16'b0000000001101100;
reg [16-1:0] bias_reg_30 = 16'b0000000000111011;
reg [16-1:0] bias_reg_31 = 16'b0000000001111101;
reg [16-1:0] bias_reg_32 = 16'b0000000001100110;
reg [16-1:0] bias_reg_33 = 16'b0000000001010000;
reg [16-1:0] bias_reg_34 = 16'b0000000001100010;
reg [16-1:0] bias_reg_35 = 16'b0000000001010011;
reg [16-1:0] bias_reg_36 = 16'b0000000001100111;
reg [16-1:0] bias_reg_37 = 16'b0000000000100100;
reg [16-1:0] bias_reg_38 = 16'b0000000001110010;
reg [16-1:0] bias_reg_39 = 16'b0000000001100101;
reg [16-1:0] bias_reg_40 = 16'b0000000001000111;
reg [16-1:0] bias_reg_41 = 16'b0000000001011011;
reg [16-1:0] bias_reg_42 = 16'b0000000001110101;
reg [16-1:0] bias_reg_43 = 16'b0000000010011001;
reg [16-1:0] bias_reg_44 = 16'b0000000000110100;
reg [16-1:0] bias_reg_45 = 16'b0000000000011111;
reg [16-1:0] bias_reg_46 = 16'b0000000010100100;
reg [16-1:0] bias_reg_47 = 16'b0000000001000011;
reg [16-1:0] bias_reg_48 = 16'b0000000001000110;
reg [16-1:0] bias_reg_49 = 16'b0000000001111101;
reg [16-1:0] bias_reg_50 = 16'b0000000000011111;
reg [16-1:0] bias_reg_51 = 16'b0000000001101110;
reg [16-1:0] bias_reg_52 = 16'b0000000001110010;
reg [16-1:0] bias_reg_53 = 16'b0000000000101111;
reg [16-1:0] bias_reg_54 = 16'b0000000000100100;
reg [16-1:0] bias_reg_55 = 16'b0000000001111100;
reg [16-1:0] bias_reg_56 = 16'b0000000000100000;
reg [16-1:0] bias_reg_57 = 16'b0000000001000100;
reg [16-1:0] bias_reg_58 = 16'b0000000001001001;
reg [16-1:0] bias_reg_59 = 16'b0000000001011011;
reg [16-1:0] bias_reg_60 = 16'b0000000001100110;
reg [16-1:0] bias_reg_61 = 16'b0000000000111011;
reg [16-1:0] bias_reg_62 = 16'b0000000001000001;
reg [16-1:0] bias_reg_63 = 16'b0000000001011100;
reg [16-1:0] bias_reg_64 = 16'b0000000001100010;
reg [16-1:0] bias_reg_65 = 16'b0000000001000000;
reg [16-1:0] bias_reg_66 = 16'b0000000000111101;
reg [16-1:0] bias_reg_67 = 16'b0000000000111111;
reg [16-1:0] bias_reg_68 = 16'b0000000001000010;
reg [16-1:0] bias_reg_69 = 16'b0000000000111111;
reg [16-1:0] bias_reg_70 = 16'b0000000001111101;
reg [16-1:0] bias_reg_71 = 16'b0000000001011101;
reg [16-1:0] bias_reg_72 = 16'b0000000000111001;
reg [16-1:0] bias_reg_73 = 16'b0000000000101010;
reg [16-1:0] bias_reg_74 = 16'b0000000000110011;
reg [16-1:0] bias_reg_75 = 16'b0000000000110000;
reg [16-1:0] bias_reg_76 = 16'b0000000000111001;
reg [16-1:0] bias_reg_77 = 16'b0000000001111100;
reg [16-1:0] bias_reg_78 = 16'b0000000001111111;
reg [16-1:0] bias_reg_79 = 16'b0000000001000000;
reg [16-1:0] bias_reg_80 = 16'b0000000001110110;
reg [16-1:0] bias_reg_81 = 16'b0000000001101100;
reg [16-1:0] bias_reg_82 = 16'b0000000000110001;
reg [16-1:0] bias_reg_83 = 16'b0000000000011100;
reg [16-1:0] bias_reg_84 = 16'b0000000010001110;
reg [16-1:0] bias_reg_85 = 16'b0000000000101010;
reg [16-1:0] bias_reg_86 = 16'b0000000000110100;
reg [16-1:0] bias_reg_87 = 16'b0000000000111101;
reg [16-1:0] bias_reg_88 = 16'b0000000001000110;
reg [16-1:0] bias_reg_89 = 16'b0000000001001010;
reg [16-1:0] bias_reg_90 = 16'b0000000010000100;
reg [16-1:0] bias_reg_91 = 16'b0000000010001000;
reg [16-1:0] bias_reg_92 = 16'b0000000010100011;
reg [16-1:0] bias_reg_93 = 16'b0000000001010100;
reg [16-1:0] bias_reg_94 = 16'b0000000001100010;
reg [16-1:0] bias_reg_95 = 16'b0000000010000110;
reg [16-1:0] bias_reg_96 = 16'b0000000001010110;
reg [16-1:0] bias_reg_97 = 16'b0000000001101000;
reg [16-1:0] bias_reg_98 = 16'b0000000001001110;
reg [16-1:0] bias_reg_99 = 16'b0000000000100011;
reg [16-1:0] bias_reg_100 = 16'b0000000001100001;
reg [16-1:0] bias_reg_101 = 16'b0000000001111111;
reg [16-1:0] bias_reg_102 = 16'b0000000001100010;
reg [16-1:0] bias_reg_103 = 16'b0000000001110111;
reg [16-1:0] bias_reg_104 = 16'b0000000000111110;
reg [16-1:0] bias_reg_105 = 16'b0000000000111010;
reg [16-1:0] bias_reg_106 = 16'b0000000001101011;
reg [16-1:0] bias_reg_107 = 16'b0000000001000010;
reg [16-1:0] bias_reg_108 = 16'b0000000000111011;
reg [16-1:0] bias_reg_109 = 16'b0000000001010100;
reg [16-1:0] bias_reg_110 = 16'b0000000001111010;
reg [16-1:0] bias_reg_111 = 16'b0000000000111100;
reg [16-1:0] bias_reg_112 = 16'b0000000000100001;
reg [16-1:0] bias_reg_113 = 16'b0000000000010100;
reg [16-1:0] bias_reg_114 = 16'b0000000010011001;
reg [16-1:0] bias_reg_115 = 16'b0000000000111111;
reg [16-1:0] bias_reg_116 = 16'b0000000001110001;
reg [16-1:0] bias_reg_117 = 16'b0000000000101000;
reg [16-1:0] bias_reg_118 = 16'b0000000001010011;
reg [16-1:0] bias_reg_119 = 16'b0000000001110110;
reg [16-1:0] bias_reg_120 = 16'b0000000000111000;
reg [16-1:0] bias_reg_121 = 16'b0000000001000011;
reg [16-1:0] bias_reg_122 = 16'b0000000001000010;
reg [16-1:0] bias_reg_123 = 16'b0000000001100010;
reg [16-1:0] bias_reg_124 = 16'b0000000001001010;
reg [16-1:0] bias_reg_125 = 16'b0000000001001100;
reg [16-1:0] bias_reg_126 = 16'b0000000010011111;
reg [16-1:0] bias_reg_127 = 16'b0000000001000011;
reg [16-1:0] bias_reg_128 = 16'b0000000010000110;
reg [16-1:0] bias_reg_129 = 16'b0000000000101110;
reg [16-1:0] bias_reg_130 = 16'b0000000000111000;
reg [16-1:0] bias_reg_131 = 16'b0000000001010101;
reg [16-1:0] bias_reg_132 = 16'b0000000001011111;
reg [16-1:0] bias_reg_133 = 16'b0000000000111110;
reg [16-1:0] bias_reg_134 = 16'b0000000001100010;
reg [16-1:0] bias_reg_135 = 16'b0000000010000000;
reg [16-1:0] bias_reg_136 = 16'b0000000000100111;
reg [16-1:0] bias_reg_137 = 16'b0000000010100111;
reg [16-1:0] bias_reg_138 = 16'b0000000001001011;
reg [16-1:0] bias_reg_139 = 16'b0000000001101111;
reg [16-1:0] bias_reg_140 = 16'b0000000001001001;
reg [16-1:0] bias_reg_141 = 16'b0000000001100000;
reg [16-1:0] bias_reg_142 = 16'b0000000001100111;
reg [16-1:0] bias_reg_143 = 16'b0000000001100110;
reg [16-1:0] bias_reg_144 = 16'b0000000010001101;
reg [16-1:0] bias_reg_145 = 16'b0000000000110111;
reg [16-1:0] bias_reg_146 = 16'b0000000001010001;
reg [16-1:0] bias_reg_147 = 16'b0000000001000010;
reg [16-1:0] bias_reg_148 = 16'b0000000010101011;
reg [16-1:0] bias_reg_149 = 16'b0000000001011101;
reg [16-1:0] bias_reg_150 = 16'b0000000010101011;
reg [16-1:0] bias_reg_151 = 16'b0000000000101101;
reg [16-1:0] bias_reg_152 = 16'b0000000001010110;
reg [16-1:0] bias_reg_153 = 16'b0000000000111100;
reg [16-1:0] bias_reg_154 = 16'b0000000010011010;
reg [16-1:0] bias_reg_155 = 16'b0000000000101010;
reg [16-1:0] bias_reg_156 = 16'b0000000001010110;
reg [16-1:0] bias_reg_157 = 16'b0000000001100011;
reg [16-1:0] bias_reg_158 = 16'b0000000001001010;
reg [16-1:0] bias_reg_159 = 16'b0000000010001100;
reg [16-1:0] bias_reg_160 = 16'b0000000001110110;
reg [16-1:0] bias_reg_161 = 16'b0000000001100000;
reg [16-1:0] bias_reg_162 = 16'b0000000001100000;
reg [16-1:0] bias_reg_163 = 16'b0000000000011101;
reg [16-1:0] bias_reg_164 = 16'b0000000001000000;
reg [16-1:0] bias_reg_165 = 16'b0000000001010110;
reg [16-1:0] bias_reg_166 = 16'b0000000010010010;
reg [16-1:0] bias_reg_167 = 16'b0000000001010110;
reg [16-1:0] bias_reg_168 = 16'b0000000000110011;
reg [16-1:0] bias_reg_169 = 16'b0000000001010110;
reg [16-1:0] bias_reg_170 = 16'b0000000001010110;
reg [16-1:0] bias_reg_171 = 16'b0000000001011101;
reg [16-1:0] bias_reg_172 = 16'b0000000001101100;
reg [16-1:0] bias_reg_173 = 16'b0000000000110011;
reg [16-1:0] bias_reg_174 = 16'b0000000000011011;
reg [16-1:0] bias_reg_175 = 16'b0000000000100010;
reg [16-1:0] bias_reg_176 = 16'b0000000001101111;
reg [16-1:0] bias_reg_177 = 16'b0000000010100010;
reg [16-1:0] bias_reg_178 = 16'b0000000001001101;
reg [16-1:0] bias_reg_179 = 16'b0000000010001100;
reg [16-1:0] bias_reg_180 = 16'b0000000010000101;
reg [16-1:0] bias_reg_181 = 16'b0000000010001110;
reg [16-1:0] bias_reg_182 = 16'b0000000001010111;
reg [16-1:0] bias_reg_183 = 16'b0000000000011101;
reg [16-1:0] bias_reg_184 = 16'b0000000001010011;
reg [16-1:0] bias_reg_185 = 16'b0000000001111101;
reg [16-1:0] bias_reg_186 = 16'b0000000001101010;
reg [16-1:0] bias_reg_187 = 16'b0000000000010101;
reg [16-1:0] bias_reg_188 = 16'b0000000001011101;
reg [16-1:0] bias_reg_189 = 16'b0000000001011111;
reg [16-1:0] bias_reg_190 = 16'b0000000000110011;
reg [16-1:0] bias_reg_191 = 16'b0000000001010110;
reg [16-1:0] bias_reg_192 = 16'b0000000000110011;
reg [16-1:0] bias_reg_193 = 16'b0000000001110111;
reg [16-1:0] bias_reg_194 = 16'b0000000001001010;
reg [16-1:0] bias_reg_195 = 16'b0000000001110010;
reg [16-1:0] bias_reg_196 = 16'b0000000010111011;
reg [16-1:0] bias_reg_197 = 16'b0000000001000111;
reg [16-1:0] bias_reg_198 = 16'b0000000010000101;
reg [16-1:0] bias_reg_199 = 16'b0000000000011001;
reg [16-1:0] bias_reg_200 = 16'b0000000000001010;
reg [16-1:0] bias_reg_201 = 16'b0000000001010101;
reg [16-1:0] bias_reg_202 = 16'b0000000001000101;
reg [16-1:0] bias_reg_203 = 16'b0000000001000001;
reg [16-1:0] bias_reg_204 = 16'b0000000001010011;
reg [16-1:0] bias_reg_205 = 16'b0000000001001111;
reg [16-1:0] bias_reg_206 = 16'b0000000001001001;
reg [16-1:0] bias_reg_207 = 16'b0000000001000010;
reg [16-1:0] bias_reg_208 = 16'b0000000010001000;
reg [16-1:0] bias_reg_209 = 16'b0000000001110100;
reg [16-1:0] bias_reg_210 = 16'b0000000010001101;
reg [16-1:0] bias_reg_211 = 16'b0000000000110001;
reg [16-1:0] bias_reg_212 = 16'b0000000001011010;
reg [16-1:0] bias_reg_213 = 16'b0000000001111011;
reg [16-1:0] bias_reg_214 = 16'b0000000000110001;
reg [16-1:0] bias_reg_215 = 16'b0000000000111110;
reg [16-1:0] bias_reg_216 = 16'b0000000010001000;
reg [16-1:0] bias_reg_217 = 16'b0000000001110101;
reg [16-1:0] bias_reg_218 = 16'b0000000000110001;
reg [16-1:0] bias_reg_219 = 16'b0000000010011010;
reg [16-1:0] bias_reg_220 = 16'b0000000001001010;
reg [16-1:0] bias_reg_221 = 16'b0000000001100001;
reg [16-1:0] bias_reg_222 = 16'b0000000000110101;
reg [16-1:0] bias_reg_223 = 16'b0000000001110010;
reg [16-1:0] bias_reg_224 = 16'b0000000001111101;
reg [16-1:0] bias_reg_225 = 16'b0000000001000011;
reg [16-1:0] bias_reg_226 = 16'b0000000001000101;
reg [16-1:0] bias_reg_227 = 16'b0000000000110000;
reg [16-1:0] bias_reg_228 = 16'b0000000001110001;
reg [16-1:0] bias_reg_229 = 16'b0000000001000101;
reg [16-1:0] bias_reg_230 = 16'b0000000001111011;
reg [16-1:0] bias_reg_231 = 16'b0000000001101100;
reg [16-1:0] bias_reg_232 = 16'b0000000001100001;
reg [16-1:0] bias_reg_233 = 16'b0000000000111111;
reg [16-1:0] bias_reg_234 = 16'b0000000000101011;
reg [16-1:0] bias_reg_235 = 16'b0000000001001011;
reg [16-1:0] bias_reg_236 = 16'b0000000000110001;
reg [16-1:0] bias_reg_237 = 16'b0000000010010101;
reg [16-1:0] bias_reg_238 = 16'b0000000000101110;
reg [16-1:0] bias_reg_239 = 16'b0000000010001010;
reg [16-1:0] bias_reg_240 = 16'b0000000001100000;
reg [16-1:0] bias_reg_241 = 16'b0000000000011100;
reg [16-1:0] bias_reg_242 = 16'b0000000001001000;
reg [16-1:0] bias_reg_243 = 16'b0000000010001111;
reg [16-1:0] bias_reg_244 = 16'b0000000000110100;
reg [16-1:0] bias_reg_245 = 16'b0000000010000000;
reg [16-1:0] bias_reg_246 = 16'b0000000001011111;
reg [16-1:0] bias_reg_247 = 16'b0000000001100101;
reg [16-1:0] bias_reg_248 = 16'b0000000001001001;
reg [16-1:0] bias_reg_249 = 16'b0000000010010010;
reg [16-1:0] bias_reg_250 = 16'b0000000001010000;
reg [16-1:0] bias_reg_251 = 16'b0000000001010010;
reg [16-1:0] bias_reg_252 = 16'b0000000001001100;
reg [16-1:0] bias_reg_253 = 16'b0000000000110101;
reg [16-1:0] bias_reg_254 = 16'b0000000000110101;
reg [16-1:0] bias_reg_255 = 16'b0000000000111001;
reg [16-1:0] bias_reg_256 = 16'b0000000000110011;
reg [16-1:0] bias_reg_257 = 16'b0000000000101101;
reg [16-1:0] bias_reg_258 = 16'b0000000001100000;
reg [16-1:0] bias_reg_259 = 16'b0000000001000001;
reg [16-1:0] bias_reg_260 = 16'b0000000010001000;
reg [16-1:0] bias_reg_261 = 16'b0000000010000001;
reg [16-1:0] bias_reg_262 = 16'b0000000001000100;
reg [16-1:0] bias_reg_263 = 16'b0000000010110010;
reg [16-1:0] bias_reg_264 = 16'b0000000010100000;
reg [16-1:0] bias_reg_265 = 16'b0000000001010010;
reg [16-1:0] bias_reg_266 = 16'b0000000000111111;
reg [16-1:0] bias_reg_267 = 16'b0000000000111111;
reg [16-1:0] bias_reg_268 = 16'b0000000000111100;
reg [16-1:0] bias_reg_269 = 16'b0000000000110101;
reg [16-1:0] bias_reg_270 = 16'b0000000001000110;
reg [16-1:0] bias_reg_271 = 16'b0000000001001101;
reg [16-1:0] bias_reg_272 = 16'b0000000001010101;
reg [16-1:0] bias_reg_273 = 16'b0000000010100011;
reg [16-1:0] bias_reg_274 = 16'b0000000010100010;
reg [16-1:0] bias_reg_275 = 16'b0000000000111011;
reg [16-1:0] bias_reg_276 = 16'b0000000001101001;
reg [16-1:0] bias_reg_277 = 16'b0000000001000111;
reg [16-1:0] bias_reg_278 = 16'b0000000010011000;
reg [16-1:0] bias_reg_279 = 16'b0000000000101101;
reg [16-1:0] bias_reg_280 = 16'b0000000001011010;
reg [16-1:0] bias_reg_281 = 16'b0000000001000010;
reg [16-1:0] bias_reg_282 = 16'b0000000001110110;
reg [16-1:0] bias_reg_283 = 16'b0000000000101110;
reg [16-1:0] bias_reg_284 = 16'b0000000000100111;
reg [16-1:0] bias_reg_285 = 16'b0000000001010101;
reg [16-1:0] bias_reg_286 = 16'b0000000001010001;
reg [16-1:0] bias_reg_287 = 16'b0000000000100110;
reg [16-1:0] bias_reg_288 = 16'b0000000000001110;
reg [16-1:0] bias_reg_289 = 16'b0000000001111110;
reg [16-1:0] bias_reg_290 = 16'b0000000010000101;
reg [16-1:0] bias_reg_291 = 16'b0000000000110110;
reg [16-1:0] bias_reg_292 = 16'b0000000001000000;
reg [16-1:0] bias_reg_293 = 16'b0000000000111101;
reg [16-1:0] bias_reg_294 = 16'b0000000001010110;
reg [16-1:0] bias_reg_295 = 16'b0000000000100001;
reg [16-1:0] bias_reg_296 = 16'b0000000001110011;
reg [16-1:0] bias_reg_297 = 16'b0000000000001111;
reg [16-1:0] bias_reg_298 = 16'b0000000001110111;
reg [16-1:0] bias_reg_299 = 16'b0000000000101101;
reg [16-1:0] bias_reg_300 = 16'b0000000001010101;
reg [16-1:0] bias_reg_301 = 16'b0000000001101001;
reg [16-1:0] bias_reg_302 = 16'b0000000001100000;
reg [16-1:0] bias_reg_303 = 16'b0000000001001101;
reg [16-1:0] bias_reg_304 = 16'b0000000001011000;
reg [16-1:0] bias_reg_305 = 16'b0000000000011110;
reg [16-1:0] bias_reg_306 = 16'b0000000001111110;
reg [16-1:0] bias_reg_307 = 16'b0000000001101000;
reg [16-1:0] bias_reg_308 = 16'b0000000001010100;
reg [16-1:0] bias_reg_309 = 16'b0000000011100100;
reg [16-1:0] bias_reg_310 = 16'b0000000000100100;
reg [16-1:0] bias_reg_311 = 16'b0000000001001100;
reg [16-1:0] bias_reg_312 = 16'b0000000001001110;
reg [16-1:0] bias_reg_313 = 16'b0000000000111110;
reg [16-1:0] bias_reg_314 = 16'b0000000010111101;
reg [16-1:0] bias_reg_315 = 16'b0000000001110100;
reg [16-1:0] bias_reg_316 = 16'b0000000001000000;
reg [16-1:0] bias_reg_317 = 16'b0000000001111001;
reg [16-1:0] bias_reg_318 = 16'b0000000001100100;
reg [16-1:0] bias_reg_319 = 16'b0000000000011010;
reg [16-1:0] bias_reg_320 = 16'b0000000001010011;
reg [16-1:0] bias_reg_321 = 16'b0000000001100110;
reg [16-1:0] bias_reg_322 = 16'b0000000000110000;
reg [16-1:0] bias_reg_323 = 16'b0000000001001101;
reg [16-1:0] bias_reg_324 = 16'b0000000001000001;
reg [16-1:0] bias_reg_325 = 16'b0000000001001110;
reg [16-1:0] bias_reg_326 = 16'b0000000001110011;
reg [16-1:0] bias_reg_327 = 16'b0000000000001101;
reg [16-1:0] bias_reg_328 = 16'b0000000001101010;
reg [16-1:0] bias_reg_329 = 16'b0000000010111111;
reg [16-1:0] bias_reg_330 = 16'b0000000001011101;
reg [16-1:0] bias_reg_331 = 16'b0000000001101101;
reg [16-1:0] bias_reg_332 = 16'b0000000001011100;
reg [16-1:0] bias_reg_333 = 16'b0000000001010100;
reg [16-1:0] bias_reg_334 = 16'b0000000000101100;
reg [16-1:0] bias_reg_335 = 16'b0000000001010100;
reg [16-1:0] bias_reg_336 = 16'b0000000001001110;
reg [16-1:0] bias_reg_337 = 16'b0000000000111101;
reg [16-1:0] bias_reg_338 = 16'b0000000000110101;
reg [16-1:0] bias_reg_339 = 16'b0000000001110010;
reg [16-1:0] bias_reg_340 = 16'b0000000000110000;
reg [16-1:0] bias_reg_341 = 16'b1000000000100110;
reg [16-1:0] bias_reg_342 = 16'b0000000001001111;
reg [16-1:0] bias_reg_343 = 16'b0000000001011011;
reg [16-1:0] bias_reg_344 = 16'b0000000001010100;
reg [16-1:0] bias_reg_345 = 16'b0000000001001011;
reg [16-1:0] bias_reg_346 = 16'b0000000001111111;
reg [16-1:0] bias_reg_347 = 16'b0000000001100000;
reg [16-1:0] bias_reg_348 = 16'b0000000001101110;
reg [16-1:0] bias_reg_349 = 16'b0000000001010000;
reg [16-1:0] bias_reg_350 = 16'b0000000010101010;
reg [16-1:0] bias_reg_351 = 16'b0000000001111000;
reg [16-1:0] bias_reg_352 = 16'b0000000000101001;
reg [16-1:0] bias_reg_353 = 16'b0000000001000000;
reg [16-1:0] bias_reg_354 = 16'b0000000001000101;
reg [16-1:0] bias_reg_355 = 16'b0000000001101001;
reg [16-1:0] bias_reg_356 = 16'b0000000001101110;
reg [16-1:0] bias_reg_357 = 16'b0000000001011101;
reg [16-1:0] bias_reg_358 = 16'b0000000001111100;
reg [16-1:0] bias_reg_359 = 16'b0000000000111001;
reg [16-1:0] bias_reg_360 = 16'b0000000001010000;
reg [16-1:0] bias_reg_361 = 16'b0000000010001010;
reg [16-1:0] bias_reg_362 = 16'b0000000000110101;
reg [16-1:0] bias_reg_363 = 16'b0000000000110000;
reg [16-1:0] bias_reg_364 = 16'b0000000001000111;
reg [16-1:0] bias_reg_365 = 16'b0000000001111110;
reg [16-1:0] bias_reg_366 = 16'b0000000001111110;
reg [16-1:0] bias_reg_367 = 16'b0000000001011010;
assign bias_mem[0] = bias_reg_0;
assign bias_mem[1] = bias_reg_1;
assign bias_mem[2] = bias_reg_2;
assign bias_mem[3] = bias_reg_3;
assign bias_mem[4] = bias_reg_4;
assign bias_mem[5] = bias_reg_5;
assign bias_mem[6] = bias_reg_6;
assign bias_mem[7] = bias_reg_7;
assign bias_mem[8] = bias_reg_8;
assign bias_mem[9] = bias_reg_9;
assign bias_mem[10] = bias_reg_10;
assign bias_mem[11] = bias_reg_11;
assign bias_mem[12] = bias_reg_12;
assign bias_mem[13] = bias_reg_13;
assign bias_mem[14] = bias_reg_14;
assign bias_mem[15] = bias_reg_15;
assign bias_mem[16] = bias_reg_16;
assign bias_mem[17] = bias_reg_17;
assign bias_mem[18] = bias_reg_18;
assign bias_mem[19] = bias_reg_19;
assign bias_mem[20] = bias_reg_20;
assign bias_mem[21] = bias_reg_21;
assign bias_mem[22] = bias_reg_22;
assign bias_mem[23] = bias_reg_23;
assign bias_mem[24] = bias_reg_24;
assign bias_mem[25] = bias_reg_25;
assign bias_mem[26] = bias_reg_26;
assign bias_mem[27] = bias_reg_27;
assign bias_mem[28] = bias_reg_28;
assign bias_mem[29] = bias_reg_29;
assign bias_mem[30] = bias_reg_30;
assign bias_mem[31] = bias_reg_31;
assign bias_mem[32] = bias_reg_32;
assign bias_mem[33] = bias_reg_33;
assign bias_mem[34] = bias_reg_34;
assign bias_mem[35] = bias_reg_35;
assign bias_mem[36] = bias_reg_36;
assign bias_mem[37] = bias_reg_37;
assign bias_mem[38] = bias_reg_38;
assign bias_mem[39] = bias_reg_39;
assign bias_mem[40] = bias_reg_40;
assign bias_mem[41] = bias_reg_41;
assign bias_mem[42] = bias_reg_42;
assign bias_mem[43] = bias_reg_43;
assign bias_mem[44] = bias_reg_44;
assign bias_mem[45] = bias_reg_45;
assign bias_mem[46] = bias_reg_46;
assign bias_mem[47] = bias_reg_47;
assign bias_mem[48] = bias_reg_48;
assign bias_mem[49] = bias_reg_49;
assign bias_mem[50] = bias_reg_50;
assign bias_mem[51] = bias_reg_51;
assign bias_mem[52] = bias_reg_52;
assign bias_mem[53] = bias_reg_53;
assign bias_mem[54] = bias_reg_54;
assign bias_mem[55] = bias_reg_55;
assign bias_mem[56] = bias_reg_56;
assign bias_mem[57] = bias_reg_57;
assign bias_mem[58] = bias_reg_58;
assign bias_mem[59] = bias_reg_59;
assign bias_mem[60] = bias_reg_60;
assign bias_mem[61] = bias_reg_61;
assign bias_mem[62] = bias_reg_62;
assign bias_mem[63] = bias_reg_63;
assign bias_mem[64] = bias_reg_64;
assign bias_mem[65] = bias_reg_65;
assign bias_mem[66] = bias_reg_66;
assign bias_mem[67] = bias_reg_67;
assign bias_mem[68] = bias_reg_68;
assign bias_mem[69] = bias_reg_69;
assign bias_mem[70] = bias_reg_70;
assign bias_mem[71] = bias_reg_71;
assign bias_mem[72] = bias_reg_72;
assign bias_mem[73] = bias_reg_73;
assign bias_mem[74] = bias_reg_74;
assign bias_mem[75] = bias_reg_75;
assign bias_mem[76] = bias_reg_76;
assign bias_mem[77] = bias_reg_77;
assign bias_mem[78] = bias_reg_78;
assign bias_mem[79] = bias_reg_79;
assign bias_mem[80] = bias_reg_80;
assign bias_mem[81] = bias_reg_81;
assign bias_mem[82] = bias_reg_82;
assign bias_mem[83] = bias_reg_83;
assign bias_mem[84] = bias_reg_84;
assign bias_mem[85] = bias_reg_85;
assign bias_mem[86] = bias_reg_86;
assign bias_mem[87] = bias_reg_87;
assign bias_mem[88] = bias_reg_88;
assign bias_mem[89] = bias_reg_89;
assign bias_mem[90] = bias_reg_90;
assign bias_mem[91] = bias_reg_91;
assign bias_mem[92] = bias_reg_92;
assign bias_mem[93] = bias_reg_93;
assign bias_mem[94] = bias_reg_94;
assign bias_mem[95] = bias_reg_95;
assign bias_mem[96] = bias_reg_96;
assign bias_mem[97] = bias_reg_97;
assign bias_mem[98] = bias_reg_98;
assign bias_mem[99] = bias_reg_99;
assign bias_mem[100] = bias_reg_100;
assign bias_mem[101] = bias_reg_101;
assign bias_mem[102] = bias_reg_102;
assign bias_mem[103] = bias_reg_103;
assign bias_mem[104] = bias_reg_104;
assign bias_mem[105] = bias_reg_105;
assign bias_mem[106] = bias_reg_106;
assign bias_mem[107] = bias_reg_107;
assign bias_mem[108] = bias_reg_108;
assign bias_mem[109] = bias_reg_109;
assign bias_mem[110] = bias_reg_110;
assign bias_mem[111] = bias_reg_111;
assign bias_mem[112] = bias_reg_112;
assign bias_mem[113] = bias_reg_113;
assign bias_mem[114] = bias_reg_114;
assign bias_mem[115] = bias_reg_115;
assign bias_mem[116] = bias_reg_116;
assign bias_mem[117] = bias_reg_117;
assign bias_mem[118] = bias_reg_118;
assign bias_mem[119] = bias_reg_119;
assign bias_mem[120] = bias_reg_120;
assign bias_mem[121] = bias_reg_121;
assign bias_mem[122] = bias_reg_122;
assign bias_mem[123] = bias_reg_123;
assign bias_mem[124] = bias_reg_124;
assign bias_mem[125] = bias_reg_125;
assign bias_mem[126] = bias_reg_126;
assign bias_mem[127] = bias_reg_127;
assign bias_mem[128] = bias_reg_128;
assign bias_mem[129] = bias_reg_129;
assign bias_mem[130] = bias_reg_130;
assign bias_mem[131] = bias_reg_131;
assign bias_mem[132] = bias_reg_132;
assign bias_mem[133] = bias_reg_133;
assign bias_mem[134] = bias_reg_134;
assign bias_mem[135] = bias_reg_135;
assign bias_mem[136] = bias_reg_136;
assign bias_mem[137] = bias_reg_137;
assign bias_mem[138] = bias_reg_138;
assign bias_mem[139] = bias_reg_139;
assign bias_mem[140] = bias_reg_140;
assign bias_mem[141] = bias_reg_141;
assign bias_mem[142] = bias_reg_142;
assign bias_mem[143] = bias_reg_143;
assign bias_mem[144] = bias_reg_144;
assign bias_mem[145] = bias_reg_145;
assign bias_mem[146] = bias_reg_146;
assign bias_mem[147] = bias_reg_147;
assign bias_mem[148] = bias_reg_148;
assign bias_mem[149] = bias_reg_149;
assign bias_mem[150] = bias_reg_150;
assign bias_mem[151] = bias_reg_151;
assign bias_mem[152] = bias_reg_152;
assign bias_mem[153] = bias_reg_153;
assign bias_mem[154] = bias_reg_154;
assign bias_mem[155] = bias_reg_155;
assign bias_mem[156] = bias_reg_156;
assign bias_mem[157] = bias_reg_157;
assign bias_mem[158] = bias_reg_158;
assign bias_mem[159] = bias_reg_159;
assign bias_mem[160] = bias_reg_160;
assign bias_mem[161] = bias_reg_161;
assign bias_mem[162] = bias_reg_162;
assign bias_mem[163] = bias_reg_163;
assign bias_mem[164] = bias_reg_164;
assign bias_mem[165] = bias_reg_165;
assign bias_mem[166] = bias_reg_166;
assign bias_mem[167] = bias_reg_167;
assign bias_mem[168] = bias_reg_168;
assign bias_mem[169] = bias_reg_169;
assign bias_mem[170] = bias_reg_170;
assign bias_mem[171] = bias_reg_171;
assign bias_mem[172] = bias_reg_172;
assign bias_mem[173] = bias_reg_173;
assign bias_mem[174] = bias_reg_174;
assign bias_mem[175] = bias_reg_175;
assign bias_mem[176] = bias_reg_176;
assign bias_mem[177] = bias_reg_177;
assign bias_mem[178] = bias_reg_178;
assign bias_mem[179] = bias_reg_179;
assign bias_mem[180] = bias_reg_180;
assign bias_mem[181] = bias_reg_181;
assign bias_mem[182] = bias_reg_182;
assign bias_mem[183] = bias_reg_183;
assign bias_mem[184] = bias_reg_184;
assign bias_mem[185] = bias_reg_185;
assign bias_mem[186] = bias_reg_186;
assign bias_mem[187] = bias_reg_187;
assign bias_mem[188] = bias_reg_188;
assign bias_mem[189] = bias_reg_189;
assign bias_mem[190] = bias_reg_190;
assign bias_mem[191] = bias_reg_191;
assign bias_mem[192] = bias_reg_192;
assign bias_mem[193] = bias_reg_193;
assign bias_mem[194] = bias_reg_194;
assign bias_mem[195] = bias_reg_195;
assign bias_mem[196] = bias_reg_196;
assign bias_mem[197] = bias_reg_197;
assign bias_mem[198] = bias_reg_198;
assign bias_mem[199] = bias_reg_199;
assign bias_mem[200] = bias_reg_200;
assign bias_mem[201] = bias_reg_201;
assign bias_mem[202] = bias_reg_202;
assign bias_mem[203] = bias_reg_203;
assign bias_mem[204] = bias_reg_204;
assign bias_mem[205] = bias_reg_205;
assign bias_mem[206] = bias_reg_206;
assign bias_mem[207] = bias_reg_207;
assign bias_mem[208] = bias_reg_208;
assign bias_mem[209] = bias_reg_209;
assign bias_mem[210] = bias_reg_210;
assign bias_mem[211] = bias_reg_211;
assign bias_mem[212] = bias_reg_212;
assign bias_mem[213] = bias_reg_213;
assign bias_mem[214] = bias_reg_214;
assign bias_mem[215] = bias_reg_215;
assign bias_mem[216] = bias_reg_216;
assign bias_mem[217] = bias_reg_217;
assign bias_mem[218] = bias_reg_218;
assign bias_mem[219] = bias_reg_219;
assign bias_mem[220] = bias_reg_220;
assign bias_mem[221] = bias_reg_221;
assign bias_mem[222] = bias_reg_222;
assign bias_mem[223] = bias_reg_223;
assign bias_mem[224] = bias_reg_224;
assign bias_mem[225] = bias_reg_225;
assign bias_mem[226] = bias_reg_226;
assign bias_mem[227] = bias_reg_227;
assign bias_mem[228] = bias_reg_228;
assign bias_mem[229] = bias_reg_229;
assign bias_mem[230] = bias_reg_230;
assign bias_mem[231] = bias_reg_231;
assign bias_mem[232] = bias_reg_232;
assign bias_mem[233] = bias_reg_233;
assign bias_mem[234] = bias_reg_234;
assign bias_mem[235] = bias_reg_235;
assign bias_mem[236] = bias_reg_236;
assign bias_mem[237] = bias_reg_237;
assign bias_mem[238] = bias_reg_238;
assign bias_mem[239] = bias_reg_239;
assign bias_mem[240] = bias_reg_240;
assign bias_mem[241] = bias_reg_241;
assign bias_mem[242] = bias_reg_242;
assign bias_mem[243] = bias_reg_243;
assign bias_mem[244] = bias_reg_244;
assign bias_mem[245] = bias_reg_245;
assign bias_mem[246] = bias_reg_246;
assign bias_mem[247] = bias_reg_247;
assign bias_mem[248] = bias_reg_248;
assign bias_mem[249] = bias_reg_249;
assign bias_mem[250] = bias_reg_250;
assign bias_mem[251] = bias_reg_251;
assign bias_mem[252] = bias_reg_252;
assign bias_mem[253] = bias_reg_253;
assign bias_mem[254] = bias_reg_254;
assign bias_mem[255] = bias_reg_255;
assign bias_mem[256] = bias_reg_256;
assign bias_mem[257] = bias_reg_257;
assign bias_mem[258] = bias_reg_258;
assign bias_mem[259] = bias_reg_259;
assign bias_mem[260] = bias_reg_260;
assign bias_mem[261] = bias_reg_261;
assign bias_mem[262] = bias_reg_262;
assign bias_mem[263] = bias_reg_263;
assign bias_mem[264] = bias_reg_264;
assign bias_mem[265] = bias_reg_265;
assign bias_mem[266] = bias_reg_266;
assign bias_mem[267] = bias_reg_267;
assign bias_mem[268] = bias_reg_268;
assign bias_mem[269] = bias_reg_269;
assign bias_mem[270] = bias_reg_270;
assign bias_mem[271] = bias_reg_271;
assign bias_mem[272] = bias_reg_272;
assign bias_mem[273] = bias_reg_273;
assign bias_mem[274] = bias_reg_274;
assign bias_mem[275] = bias_reg_275;
assign bias_mem[276] = bias_reg_276;
assign bias_mem[277] = bias_reg_277;
assign bias_mem[278] = bias_reg_278;
assign bias_mem[279] = bias_reg_279;
assign bias_mem[280] = bias_reg_280;
assign bias_mem[281] = bias_reg_281;
assign bias_mem[282] = bias_reg_282;
assign bias_mem[283] = bias_reg_283;
assign bias_mem[284] = bias_reg_284;
assign bias_mem[285] = bias_reg_285;
assign bias_mem[286] = bias_reg_286;
assign bias_mem[287] = bias_reg_287;
assign bias_mem[288] = bias_reg_288;
assign bias_mem[289] = bias_reg_289;
assign bias_mem[290] = bias_reg_290;
assign bias_mem[291] = bias_reg_291;
assign bias_mem[292] = bias_reg_292;
assign bias_mem[293] = bias_reg_293;
assign bias_mem[294] = bias_reg_294;
assign bias_mem[295] = bias_reg_295;
assign bias_mem[296] = bias_reg_296;
assign bias_mem[297] = bias_reg_297;
assign bias_mem[298] = bias_reg_298;
assign bias_mem[299] = bias_reg_299;
assign bias_mem[300] = bias_reg_300;
assign bias_mem[301] = bias_reg_301;
assign bias_mem[302] = bias_reg_302;
assign bias_mem[303] = bias_reg_303;
assign bias_mem[304] = bias_reg_304;
assign bias_mem[305] = bias_reg_305;
assign bias_mem[306] = bias_reg_306;
assign bias_mem[307] = bias_reg_307;
assign bias_mem[308] = bias_reg_308;
assign bias_mem[309] = bias_reg_309;
assign bias_mem[310] = bias_reg_310;
assign bias_mem[311] = bias_reg_311;
assign bias_mem[312] = bias_reg_312;
assign bias_mem[313] = bias_reg_313;
assign bias_mem[314] = bias_reg_314;
assign bias_mem[315] = bias_reg_315;
assign bias_mem[316] = bias_reg_316;
assign bias_mem[317] = bias_reg_317;
assign bias_mem[318] = bias_reg_318;
assign bias_mem[319] = bias_reg_319;
assign bias_mem[320] = bias_reg_320;
assign bias_mem[321] = bias_reg_321;
assign bias_mem[322] = bias_reg_322;
assign bias_mem[323] = bias_reg_323;
assign bias_mem[324] = bias_reg_324;
assign bias_mem[325] = bias_reg_325;
assign bias_mem[326] = bias_reg_326;
assign bias_mem[327] = bias_reg_327;
assign bias_mem[328] = bias_reg_328;
assign bias_mem[329] = bias_reg_329;
assign bias_mem[330] = bias_reg_330;
assign bias_mem[331] = bias_reg_331;
assign bias_mem[332] = bias_reg_332;
assign bias_mem[333] = bias_reg_333;
assign bias_mem[334] = bias_reg_334;
assign bias_mem[335] = bias_reg_335;
assign bias_mem[336] = bias_reg_336;
assign bias_mem[337] = bias_reg_337;
assign bias_mem[338] = bias_reg_338;
assign bias_mem[339] = bias_reg_339;
assign bias_mem[340] = bias_reg_340;
assign bias_mem[341] = bias_reg_341;
assign bias_mem[342] = bias_reg_342;
assign bias_mem[343] = bias_reg_343;
assign bias_mem[344] = bias_reg_344;
assign bias_mem[345] = bias_reg_345;
assign bias_mem[346] = bias_reg_346;
assign bias_mem[347] = bias_reg_347;
assign bias_mem[348] = bias_reg_348;
assign bias_mem[349] = bias_reg_349;
assign bias_mem[350] = bias_reg_350;
assign bias_mem[351] = bias_reg_351;
assign bias_mem[352] = bias_reg_352;
assign bias_mem[353] = bias_reg_353;
assign bias_mem[354] = bias_reg_354;
assign bias_mem[355] = bias_reg_355;
assign bias_mem[356] = bias_reg_356;
assign bias_mem[357] = bias_reg_357;
assign bias_mem[358] = bias_reg_358;
assign bias_mem[359] = bias_reg_359;
assign bias_mem[360] = bias_reg_360;
assign bias_mem[361] = bias_reg_361;
assign bias_mem[362] = bias_reg_362;
assign bias_mem[363] = bias_reg_363;
assign bias_mem[364] = bias_reg_364;
assign bias_mem[365] = bias_reg_365;
assign bias_mem[366] = bias_reg_366;
assign bias_mem[367] = bias_reg_367;
endmodule
